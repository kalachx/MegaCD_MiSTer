module composite_pal
(
    input clk, 
    input [11:0] index,
    output reg [23:0] out
);

always @ (posedge clk)
    case (index)
        12'd0000: out <= 24'h000000;
        12'd0001: out <= 24'h00000e;
        12'd0002: out <= 24'h00001b;
        12'd0003: out <= 24'h00012c;
        12'd0004: out <= 24'h01023d;
        12'd0005: out <= 24'h00014a;
        12'd0006: out <= 24'h000058;
        12'd0007: out <= 24'h00026a;
        12'd0008: out <= 24'h01047b;
        12'd0009: out <= 24'h000288;
        12'd0010: out <= 24'h000095;
        12'd0011: out <= 24'h0102a6;
        12'd0012: out <= 24'h0205b8;
        12'd0013: out <= 24'h0104c6;
        12'd0014: out <= 24'h0002d3;
        12'd0015: out <= 24'h0002d3;
        12'd0016: out <= 24'h041201;
        12'd0017: out <= 24'h02110e;
        12'd0018: out <= 24'h02111c;
        12'd0019: out <= 24'h04142e;
        12'd0020: out <= 24'h05143e;
        12'd0021: out <= 24'h04134c;
        12'd0022: out <= 24'h031259;
        12'd0023: out <= 24'h05146a;
        12'd0024: out <= 24'h06167c;
        12'd0025: out <= 24'h04148a;
        12'd0026: out <= 24'h031296;
        12'd0027: out <= 24'h0615a8;
        12'd0028: out <= 24'h0618b9;
        12'd0029: out <= 24'h0416c6;
        12'd0030: out <= 24'h0414d4;
        12'd0031: out <= 24'h0414d4;
        12'd0032: out <= 24'h092502;
        12'd0033: out <= 24'h072410;
        12'd0034: out <= 24'h05221d;
        12'd0035: out <= 24'h07242e;
        12'd0036: out <= 24'h092740;
        12'd0037: out <= 24'h08264d;
        12'd0038: out <= 24'h06245a;
        12'd0039: out <= 24'h08266c;
        12'd0040: out <= 24'h0a297d;
        12'd0041: out <= 24'h08278a;
        12'd0042: out <= 24'h062598;
        12'd0043: out <= 24'h0828a9;
        12'd0044: out <= 24'h0b2aba;
        12'd0045: out <= 24'h0928c8;
        12'd0046: out <= 24'h0727d5;
        12'd0047: out <= 24'h0727d5;
        12'd0048: out <= 24'h093401;
        12'd0049: out <= 24'h0c3610;
        12'd0050: out <= 24'h0a341e;
        12'd0051: out <= 24'h08332c;
        12'd0052: out <= 24'h0a363d;
        12'd0053: out <= 24'h0c384e;
        12'd0054: out <= 24'h0a365b;
        12'd0055: out <= 24'h083568;
        12'd0056: out <= 24'h0a387a;
        12'd0057: out <= 24'h0c3a8c;
        12'd0058: out <= 24'h0a3899;
        12'd0059: out <= 24'h0836a6;
        12'd0060: out <= 24'h0b38b7;
        12'd0061: out <= 24'h0e3bc8;
        12'd0062: out <= 24'h0c3ad6;
        12'd0063: out <= 24'h0c3ad6;
        12'd0064: out <= 24'h094200;
        12'd0065: out <= 24'h0c4410;
        12'd0066: out <= 24'h0e471f;
        12'd0067: out <= 24'h0c462c;
        12'd0068: out <= 24'h0a443a;
        12'd0069: out <= 24'h0c464b;
        12'd0070: out <= 24'h0e495c;
        12'd0071: out <= 24'h0c486a;
        12'd0072: out <= 24'h0a4677;
        12'd0073: out <= 24'h0c4888;
        12'd0074: out <= 24'h0f4b9a;
        12'd0075: out <= 24'h0d49a7;
        12'd0076: out <= 24'h0b47b4;
        12'd0077: out <= 24'h0e4ac6;
        12'd0078: out <= 24'h104cd7;
        12'd0079: out <= 24'h104cd7;
        12'd0080: out <= 24'h0e5400;
        12'd0081: out <= 24'h0c530c;
        12'd0082: out <= 24'h0e561c;
        12'd0083: out <= 24'h10582e;
        12'd0084: out <= 24'h0e563b;
        12'd0085: out <= 24'h0c5548;
        12'd0086: out <= 24'h0e5859;
        12'd0087: out <= 24'h105a6a;
        12'd0088: out <= 24'h0e5878;
        12'd0089: out <= 24'h0c5786;
        12'd0090: out <= 24'h0f5a97;
        12'd0091: out <= 24'h125ca8;
        12'd0092: out <= 24'h105ab6;
        12'd0093: out <= 24'h0e58c2;
        12'd0094: out <= 24'h105ad4;
        12'd0095: out <= 24'h105ad4;
        12'd0096: out <= 24'h126700;
        12'd0097: out <= 24'h10660c;
        12'd0098: out <= 24'h0e6419;
        12'd0099: out <= 24'h10662a;
        12'd0100: out <= 24'h12693c;
        12'd0101: out <= 24'h106849;
        12'd0102: out <= 24'h0f6656;
        12'd0103: out <= 24'h116868;
        12'd0104: out <= 24'h136b79;
        12'd0105: out <= 24'h116a86;
        12'd0106: out <= 24'h0f6894;
        12'd0107: out <= 24'h126aa6;
        12'd0108: out <= 24'h146db7;
        12'd0109: out <= 24'h126bc4;
        12'd0110: out <= 24'h1069d1;
        12'd0111: out <= 24'h1069d1;
        12'd0112: out <= 24'h127600;
        12'd0113: out <= 24'h14780e;
        12'd0114: out <= 24'h12761a;
        12'd0115: out <= 24'h107528;
        12'd0116: out <= 24'h127839;
        12'd0117: out <= 24'h147a4a;
        12'd0118: out <= 24'h137858;
        12'd0119: out <= 24'h127764;
        12'd0120: out <= 24'h147a76;
        12'd0121: out <= 24'h167c88;
        12'd0122: out <= 24'h147a95;
        12'd0123: out <= 24'h1279a2;
        12'd0124: out <= 24'h147cb4;
        12'd0125: out <= 24'h167ec5;
        12'd0126: out <= 24'h147cd2;
        12'd0127: out <= 24'h147cd2;
        12'd0128: out <= 24'h128400;
        12'd0129: out <= 24'h14860e;
        12'd0130: out <= 24'h17891b;
        12'd0131: out <= 24'h158828;
        12'd0132: out <= 24'h138636;
        12'd0133: out <= 24'h158848;
        12'd0134: out <= 24'h178b59;
        12'd0135: out <= 24'h168a66;
        12'd0136: out <= 24'h148873;
        12'd0137: out <= 24'h168a84;
        12'd0138: out <= 24'h188d96;
        12'd0139: out <= 24'h168ca4;
        12'd0140: out <= 24'h148ab1;
        12'd0141: out <= 24'h168cc2;
        12'd0142: out <= 24'h198fd3;
        12'd0143: out <= 24'h198fd3;
        12'd0144: out <= 24'h169600;
        12'd0145: out <= 24'h18990f;
        12'd0146: out <= 24'h1b9c1c;
        12'd0147: out <= 24'h1a9a2a;
        12'd0148: out <= 24'h189837;
        12'd0149: out <= 24'h1a9b48;
        12'd0150: out <= 24'h1c9e5a;
        12'd0151: out <= 24'h1a9c68;
        12'd0152: out <= 24'h189a74;
        12'd0153: out <= 24'h1a9d86;
        12'd0154: out <= 24'h1ca097;
        12'd0155: out <= 24'h1a9ea4;
        12'd0156: out <= 24'h189cb2;
        12'd0157: out <= 24'h169abf;
        12'd0158: out <= 24'h199dd0;
        12'd0159: out <= 24'h199dd0;
        12'd0160: out <= 24'h1ba900;
        12'd0161: out <= 24'h1dac0f;
        12'd0162: out <= 24'h1fae1e;
        12'd0163: out <= 24'h1eac2b;
        12'd0164: out <= 24'h1cab38;
        12'd0165: out <= 24'h1eae4a;
        12'd0166: out <= 24'h20b05b;
        12'd0167: out <= 24'h1eae68;
        12'd0168: out <= 24'h1cad76;
        12'd0169: out <= 24'h1eb087;
        12'd0170: out <= 24'h21b298;
        12'd0171: out <= 24'h1fb0a6;
        12'd0172: out <= 24'h1dafb3;
        12'd0173: out <= 24'h1badc0;
        12'd0174: out <= 24'h19abcd;
        12'd0175: out <= 24'h19abcd;
        12'd0176: out <= 24'h20bc00;
        12'd0177: out <= 24'h1eba0c;
        12'd0178: out <= 24'h20bc1b;
        12'd0179: out <= 24'h22bf2c;
        12'd0180: out <= 24'h20be39;
        12'd0181: out <= 24'h1ebc46;
        12'd0182: out <= 24'h20be58;
        12'd0183: out <= 24'h22c16a;
        12'd0184: out <= 24'h20c077;
        12'd0185: out <= 24'h1ebe84;
        12'd0186: out <= 24'h21c095;
        12'd0187: out <= 24'h24c3a6;
        12'd0188: out <= 24'h22c2b4;
        12'd0189: out <= 24'h20c0c2;
        12'd0190: out <= 24'h1ebece;
        12'd0191: out <= 24'h1ebece;
        12'd0192: out <= 24'h24cf00;
        12'd0193: out <= 24'h22cd0c;
        12'd0194: out <= 24'h20cb18;
        12'd0195: out <= 24'h22ce29;
        12'd0196: out <= 24'h24d03a;
        12'd0197: out <= 24'h22ce48;
        12'd0198: out <= 24'h21cd55;
        12'd0199: out <= 24'h23d066;
        12'd0200: out <= 24'h25d278;
        12'd0201: out <= 24'h23d085;
        12'd0202: out <= 24'h21cf92;
        12'd0203: out <= 24'h24d2a4;
        12'd0204: out <= 24'h26d4b5;
        12'd0205: out <= 24'h24d2c2;
        12'd0206: out <= 24'h22d1d0;
        12'd0207: out <= 24'h22d1d0;
        12'd0208: out <= 24'h24de00;
        12'd0209: out <= 24'h26e00d;
        12'd0210: out <= 24'h24de19;
        12'd0211: out <= 24'h22dc26;
        12'd0212: out <= 24'h24de37;
        12'd0213: out <= 24'h26e148;
        12'd0214: out <= 24'h25e056;
        12'd0215: out <= 24'h23de64;
        12'd0216: out <= 24'h25e075;
        12'd0217: out <= 24'h28e386;
        12'd0218: out <= 24'h26e294;
        12'd0219: out <= 24'h24e0a0;
        12'd0220: out <= 24'h26e2b2;
        12'd0221: out <= 24'h28e5c4;
        12'd0222: out <= 24'h26e4d1;
        12'd0223: out <= 24'h26e4d1;
        12'd0224: out <= 24'h24ec00;
        12'd0225: out <= 24'h26ee0d;
        12'd0226: out <= 24'h29f11a;
        12'd0227: out <= 24'h27ef27;
        12'd0228: out <= 24'h25ed34;
        12'd0229: out <= 24'h27f046;
        12'd0230: out <= 24'h29f257;
        12'd0231: out <= 24'h27f064;
        12'd0232: out <= 24'h25ef72;
        12'd0233: out <= 24'h28f284;
        12'd0234: out <= 24'h2af495;
        12'd0235: out <= 24'h28f2a2;
        12'd0236: out <= 24'h26f1af;
        12'd0237: out <= 24'h28f4c0;
        12'd0238: out <= 24'h2bf6d2;
        12'd0239: out <= 24'h2bf6d2;
        12'd0240: out <= 24'h24ec00;
        12'd0241: out <= 24'h26ee0d;
        12'd0242: out <= 24'h29f11a;
        12'd0243: out <= 24'h27ef27;
        12'd0244: out <= 24'h25ed34;
        12'd0245: out <= 24'h27f046;
        12'd0246: out <= 24'h29f257;
        12'd0247: out <= 24'h27f064;
        12'd0248: out <= 24'h25ef72;
        12'd0249: out <= 24'h28f284;
        12'd0250: out <= 24'h2af495;
        12'd0251: out <= 24'h28f2a2;
        12'd0252: out <= 24'h26f1af;
        12'd0253: out <= 24'h28f4c0;
        12'd0254: out <= 24'h2bf6d2;
        12'd0255: out <= 24'h2bf6d2;
        12'd0256: out <= 24'h0e0002;
        12'd0257: out <= 24'h100214;
        12'd0258: out <= 24'h100221;
        12'd0259: out <= 24'h0e002e;
        12'd0260: out <= 24'h0f023f;
        12'd0261: out <= 24'h110450;
        12'd0262: out <= 24'h10035e;
        12'd0263: out <= 24'h0e016c;
        12'd0264: out <= 24'h0f037d;
        12'd0265: out <= 24'h12068e;
        12'd0266: out <= 24'h11049c;
        12'd0267: out <= 24'h0f02a8;
        12'd0268: out <= 24'h1004ba;
        12'd0269: out <= 24'h1207cc;
        12'd0270: out <= 24'h1106d9;
        12'd0271: out <= 24'h1106d9;
        12'd0272: out <= 24'h121203;
        12'd0273: out <= 24'h101010;
        12'd0274: out <= 24'h10101e;
        12'd0275: out <= 24'h121330;
        12'd0276: out <= 24'h131440;
        12'd0277: out <= 24'h12124e;
        12'd0278: out <= 24'h11125b;
        12'd0279: out <= 24'h13146c;
        12'd0280: out <= 24'h14167e;
        12'd0281: out <= 24'h12148c;
        12'd0282: out <= 24'h111298;
        12'd0283: out <= 24'h1414aa;
        12'd0284: out <= 24'h1417bb;
        12'd0285: out <= 24'h1216c8;
        12'd0286: out <= 24'h1214d6;
        12'd0287: out <= 24'h1214d6;
        12'd0288: out <= 24'h172404;
        12'd0289: out <= 24'h152312;
        12'd0290: out <= 24'h13221f;
        12'd0291: out <= 24'h152430;
        12'd0292: out <= 24'h172642;
        12'd0293: out <= 24'h16254f;
        12'd0294: out <= 24'h14245c;
        12'd0295: out <= 24'h16266e;
        12'd0296: out <= 24'h18287f;
        12'd0297: out <= 24'h16268c;
        12'd0298: out <= 24'h14249a;
        12'd0299: out <= 24'h1627ab;
        12'd0300: out <= 24'h192abc;
        12'd0301: out <= 24'h1728ca;
        12'd0302: out <= 24'h1526d7;
        12'd0303: out <= 24'h1526d7;
        12'd0304: out <= 24'h1b3706;
        12'd0305: out <= 24'h1a3612;
        12'd0306: out <= 24'h183420;
        12'd0307: out <= 24'h1a3632;
        12'd0308: out <= 24'h1c3943;
        12'd0309: out <= 24'h1a3850;
        12'd0310: out <= 24'h18365e;
        12'd0311: out <= 24'h1a386e;
        12'd0312: out <= 24'h1c3b80;
        12'd0313: out <= 24'h1a3a8e;
        12'd0314: out <= 24'h18389b;
        12'd0315: out <= 24'h1636a8;
        12'd0316: out <= 24'h1938b9;
        12'd0317: out <= 24'h1c3aca;
        12'd0318: out <= 24'h1a39d8;
        12'd0319: out <= 24'h1a39d8;
        12'd0320: out <= 24'h1b4604;
        12'd0321: out <= 24'h1a4412;
        12'd0322: out <= 24'h1c4621;
        12'd0323: out <= 24'h1e4932;
        12'd0324: out <= 24'h1c4840;
        12'd0325: out <= 24'h1a464e;
        12'd0326: out <= 24'h1c485e;
        12'd0327: out <= 24'h1e4b70;
        12'd0328: out <= 24'h1c4a7d;
        12'd0329: out <= 24'h1a488a;
        12'd0330: out <= 24'h1d4a9c;
        12'd0331: out <= 24'h1b48a9;
        12'd0332: out <= 24'h1946b6;
        12'd0333: out <= 24'h1c49c8;
        12'd0334: out <= 24'h1e4cd9;
        12'd0335: out <= 24'h1e4cd9;
        12'd0336: out <= 24'h1c5402;
        12'd0337: out <= 24'h1e5612;
        12'd0338: out <= 24'h205922;
        12'd0339: out <= 24'h1e5830;
        12'd0340: out <= 24'h1c563d;
        12'd0341: out <= 24'h1e584e;
        12'd0342: out <= 24'h205b60;
        12'd0343: out <= 24'h1e5a6c;
        12'd0344: out <= 24'h1c587a;
        12'd0345: out <= 24'h1f5a8c;
        12'd0346: out <= 24'h225d9d;
        12'd0347: out <= 24'h205caa;
        12'd0348: out <= 24'h1e5ab8;
        12'd0349: out <= 24'h205cc8;
        12'd0350: out <= 24'h225eda;
        12'd0351: out <= 24'h225eda;
        12'd0352: out <= 24'h206602;
        12'd0353: out <= 24'h226912;
        12'd0354: out <= 24'h20681f;
        12'd0355: out <= 24'h1e662c;
        12'd0356: out <= 24'h20683e;
        12'd0357: out <= 24'h226b50;
        12'd0358: out <= 24'h216a5c;
        12'd0359: out <= 24'h1f686a;
        12'd0360: out <= 24'h216a7b;
        12'd0361: out <= 24'h246d8c;
        12'd0362: out <= 24'h226c9a;
        12'd0363: out <= 24'h206aa8;
        12'd0364: out <= 24'h226cb9;
        12'd0365: out <= 24'h246fca;
        12'd0366: out <= 24'h226dd7;
        12'd0367: out <= 24'h226dd7;
        12'd0368: out <= 24'h247902;
        12'd0369: out <= 24'h227810;
        12'd0370: out <= 24'h20761c;
        12'd0371: out <= 24'h22782e;
        12'd0372: out <= 24'h247b3f;
        12'd0373: out <= 24'h227a4c;
        12'd0374: out <= 24'h21785a;
        12'd0375: out <= 24'h247a6b;
        12'd0376: out <= 24'h267d7c;
        12'd0377: out <= 24'h247c8a;
        12'd0378: out <= 24'h227a97;
        12'd0379: out <= 24'h247ca8;
        12'd0380: out <= 24'h267fba;
        12'd0381: out <= 24'h247dc7;
        12'd0382: out <= 24'h227bd4;
        12'd0383: out <= 24'h227bd4;
        12'd0384: out <= 24'h248802;
        12'd0385: out <= 24'h228610;
        12'd0386: out <= 24'h25881d;
        12'd0387: out <= 24'h278b2e;
        12'd0388: out <= 24'h258a3c;
        12'd0389: out <= 24'h23884a;
        12'd0390: out <= 24'h258a5b;
        12'd0391: out <= 24'h288d6c;
        12'd0392: out <= 24'h268c7a;
        12'd0393: out <= 24'h248a86;
        12'd0394: out <= 24'h268c98;
        12'd0395: out <= 24'h288faa;
        12'd0396: out <= 24'h268eb7;
        12'd0397: out <= 24'h248cc4;
        12'd0398: out <= 24'h278ed5;
        12'd0399: out <= 24'h278ed5;
        12'd0400: out <= 24'h249600;
        12'd0401: out <= 24'h269811;
        12'd0402: out <= 24'h299b1e;
        12'd0403: out <= 24'h289a2c;
        12'd0404: out <= 24'h269839;
        12'd0405: out <= 24'h289a4a;
        12'd0406: out <= 24'h2a9d5c;
        12'd0407: out <= 24'h289c6a;
        12'd0408: out <= 24'h269a76;
        12'd0409: out <= 24'h289c88;
        12'd0410: out <= 24'h2a9f99;
        12'd0411: out <= 24'h289ea6;
        12'd0412: out <= 24'h269cb4;
        12'd0413: out <= 24'h289ec6;
        12'd0414: out <= 24'h2ba1d6;
        12'd0415: out <= 24'h2ba1d6;
        12'd0416: out <= 24'h29a800;
        12'd0417: out <= 24'h2bab11;
        12'd0418: out <= 24'h2dae20;
        12'd0419: out <= 24'h2cac2d;
        12'd0420: out <= 24'h2aaa3a;
        12'd0421: out <= 24'h2cad4c;
        12'd0422: out <= 24'h2eb05d;
        12'd0423: out <= 24'h2cae6a;
        12'd0424: out <= 24'h2aac78;
        12'd0425: out <= 24'h2caf89;
        12'd0426: out <= 24'h2fb29a;
        12'd0427: out <= 24'h2db0a8;
        12'd0428: out <= 24'h2baeb5;
        12'd0429: out <= 24'h2db1c6;
        12'd0430: out <= 24'h2bafd4;
        12'd0431: out <= 24'h2bafd4;
        12'd0432: out <= 24'h2ebc00;
        12'd0433: out <= 24'h2cba0e;
        12'd0434: out <= 24'h2ebc1d;
        12'd0435: out <= 24'h30be2e;
        12'd0436: out <= 24'h2ebd3c;
        12'd0437: out <= 24'h2cbc48;
        12'd0438: out <= 24'h2ebe5a;
        12'd0439: out <= 24'h30c06c;
        12'd0440: out <= 24'h2ebf79;
        12'd0441: out <= 24'h2cbe86;
        12'd0442: out <= 24'h2fc097;
        12'd0443: out <= 24'h32c2a8;
        12'd0444: out <= 24'h30c1b6;
        12'd0445: out <= 24'h2ec0c4;
        12'd0446: out <= 24'h2cbed0;
        12'd0447: out <= 24'h2cbed0;
        12'd0448: out <= 24'h32ce00;
        12'd0449: out <= 24'h30cc0e;
        12'd0450: out <= 24'h2eca1a;
        12'd0451: out <= 24'h30cd2c;
        12'd0452: out <= 24'h32d03c;
        12'd0453: out <= 24'h30ce4a;
        12'd0454: out <= 24'h2fcc57;
        12'd0455: out <= 24'h31cf68;
        12'd0456: out <= 24'h33d27a;
        12'd0457: out <= 24'h31d087;
        12'd0458: out <= 24'h2fce94;
        12'd0459: out <= 24'h32d1a6;
        12'd0460: out <= 24'h34d4b7;
        12'd0461: out <= 24'h32d2c4;
        12'd0462: out <= 24'h30d0d2;
        12'd0463: out <= 24'h30d0d2;
        12'd0464: out <= 24'h36e102;
        12'd0465: out <= 24'h34e00f;
        12'd0466: out <= 24'h32de1b;
        12'd0467: out <= 24'h34e02c;
        12'd0468: out <= 24'h36e23e;
        12'd0469: out <= 24'h34e04a;
        12'd0470: out <= 24'h33df58;
        12'd0471: out <= 24'h36e26a;
        12'd0472: out <= 24'h38e47b;
        12'd0473: out <= 24'h36e288;
        12'd0474: out <= 24'h34e196;
        12'd0475: out <= 24'h36e4a6;
        12'd0476: out <= 24'h38e6b8;
        12'd0477: out <= 24'h36e4c6;
        12'd0478: out <= 24'h34e3d3;
        12'd0479: out <= 24'h34e3d3;
        12'd0480: out <= 24'h36f002;
        12'd0481: out <= 24'h34ee0f;
        12'd0482: out <= 24'h37f01c;
        12'd0483: out <= 24'h39f32e;
        12'd0484: out <= 24'h37f13a;
        12'd0485: out <= 24'h35ef48;
        12'd0486: out <= 24'h37f259;
        12'd0487: out <= 24'h3af46a;
        12'd0488: out <= 24'h38f278;
        12'd0489: out <= 24'h36f186;
        12'd0490: out <= 24'h38f497;
        12'd0491: out <= 24'h3af6a8;
        12'd0492: out <= 24'h38f4b5;
        12'd0493: out <= 24'h36f3c2;
        12'd0494: out <= 24'h39f6d4;
        12'd0495: out <= 24'h39f6d4;
        12'd0496: out <= 24'h36f002;
        12'd0497: out <= 24'h34ee0f;
        12'd0498: out <= 24'h37f01c;
        12'd0499: out <= 24'h39f32e;
        12'd0500: out <= 24'h37f13a;
        12'd0501: out <= 24'h35ef48;
        12'd0502: out <= 24'h37f259;
        12'd0503: out <= 24'h3af46a;
        12'd0504: out <= 24'h38f278;
        12'd0505: out <= 24'h36f186;
        12'd0506: out <= 24'h38f497;
        12'd0507: out <= 24'h3af6a8;
        12'd0508: out <= 24'h38f4b5;
        12'd0509: out <= 24'h36f3c2;
        12'd0510: out <= 24'h39f6d4;
        12'd0511: out <= 24'h39f6d4;
        12'd0512: out <= 24'h1c0004;
        12'd0513: out <= 24'h1e0216;
        12'd0514: out <= 24'h200427;
        12'd0515: out <= 24'h1e0234;
        12'd0516: out <= 24'h1d0141;
        12'd0517: out <= 24'h1f0452;
        12'd0518: out <= 24'h210664;
        12'd0519: out <= 24'h1f0472;
        12'd0520: out <= 24'h1d027f;
        12'd0521: out <= 24'h200490;
        12'd0522: out <= 24'h2207a2;
        12'd0523: out <= 24'h2006af;
        12'd0524: out <= 24'h1e04bc;
        12'd0525: out <= 24'h2006ce;
        12'd0526: out <= 24'h2209df;
        12'd0527: out <= 24'h2209df;
        12'd0528: out <= 24'h201205;
        12'd0529: out <= 24'h1e1012;
        12'd0530: out <= 24'h201224;
        12'd0531: out <= 24'h221536;
        12'd0532: out <= 24'h211442;
        12'd0533: out <= 24'h201250;
        12'd0534: out <= 24'h221461;
        12'd0535: out <= 24'h241772;
        12'd0536: out <= 24'h221580;
        12'd0537: out <= 24'h20138e;
        12'd0538: out <= 24'h22169f;
        12'd0539: out <= 24'h2418b0;
        12'd0540: out <= 24'h2216bd;
        12'd0541: out <= 24'h2015ca;
        12'd0542: out <= 24'h2218dc;
        12'd0543: out <= 24'h2218dc;
        12'd0544: out <= 24'h252406;
        12'd0545: out <= 24'h232214;
        12'd0546: out <= 24'h212121;
        12'd0547: out <= 24'h232432;
        12'd0548: out <= 24'h252644;
        12'd0549: out <= 24'h242451;
        12'd0550: out <= 24'h22235e;
        12'd0551: out <= 24'h242670;
        12'd0552: out <= 24'h262881;
        12'd0553: out <= 24'h24268e;
        12'd0554: out <= 24'h22249c;
        12'd0555: out <= 24'h2426ad;
        12'd0556: out <= 24'h2729be;
        12'd0557: out <= 24'h2528cc;
        12'd0558: out <= 24'h2326d9;
        12'd0559: out <= 24'h2326d9;
        12'd0560: out <= 24'h293608;
        12'd0561: out <= 24'h283514;
        12'd0562: out <= 24'h263422;
        12'd0563: out <= 24'h283634;
        12'd0564: out <= 24'h2a3845;
        12'd0565: out <= 24'h283752;
        12'd0566: out <= 24'h263660;
        12'd0567: out <= 24'h283870;
        12'd0568: out <= 24'h2a3a82;
        12'd0569: out <= 24'h283990;
        12'd0570: out <= 24'h26379d;
        12'd0571: out <= 24'h2435aa;
        12'd0572: out <= 24'h2738bb;
        12'd0573: out <= 24'h2a3acc;
        12'd0574: out <= 24'h2838da;
        12'd0575: out <= 24'h2838da;
        12'd0576: out <= 24'h2d4909;
        12'd0577: out <= 24'h2c4816;
        12'd0578: out <= 24'h2a4623;
        12'd0579: out <= 24'h2c4834;
        12'd0580: out <= 24'h2e4b46;
        12'd0581: out <= 24'h2c4a54;
        12'd0582: out <= 24'h2a4861;
        12'd0583: out <= 24'h2c4a72;
        12'd0584: out <= 24'h2f4d83;
        12'd0585: out <= 24'h2d4c90;
        12'd0586: out <= 24'h2b4a9e;
        12'd0587: out <= 24'h2948ab;
        12'd0588: out <= 24'h2746b8;
        12'd0589: out <= 24'h2a48ca;
        12'd0590: out <= 24'h2c4bdb;
        12'd0591: out <= 24'h2c4bdb;
        12'd0592: out <= 24'h2e5806;
        12'd0593: out <= 24'h305a17;
        12'd0594: out <= 24'h2e5824;
        12'd0595: out <= 24'h2c5732;
        12'd0596: out <= 24'h2e5a43;
        12'd0597: out <= 24'h305c54;
        12'd0598: out <= 24'h2e5a62;
        12'd0599: out <= 24'h2c596f;
        12'd0600: out <= 24'h2f5c80;
        12'd0601: out <= 24'h325e92;
        12'd0602: out <= 24'h305c9f;
        12'd0603: out <= 24'h2e5bac;
        12'd0604: out <= 24'h2c59ba;
        12'd0605: out <= 24'h2e5cca;
        12'd0606: out <= 24'h305edc;
        12'd0607: out <= 24'h305edc;
        12'd0608: out <= 24'h2e6603;
        12'd0609: out <= 24'h306814;
        12'd0610: out <= 24'h326b25;
        12'd0611: out <= 24'h306a32;
        12'd0612: out <= 24'h2e6840;
        12'd0613: out <= 24'h306a52;
        12'd0614: out <= 24'h336d63;
        12'd0615: out <= 24'h316c70;
        12'd0616: out <= 24'h2f6a7d;
        12'd0617: out <= 24'h326c8e;
        12'd0618: out <= 24'h346fa0;
        12'd0619: out <= 24'h326eae;
        12'd0620: out <= 24'h306cbb;
        12'd0621: out <= 24'h326ecc;
        12'd0622: out <= 24'h3471dd;
        12'd0623: out <= 24'h3471dd;
        12'd0624: out <= 24'h327804;
        12'd0625: out <= 24'h307711;
        12'd0626: out <= 24'h327a22;
        12'd0627: out <= 24'h347c34;
        12'd0628: out <= 24'h327a41;
        12'd0629: out <= 24'h30794e;
        12'd0630: out <= 24'h337c60;
        12'd0631: out <= 24'h367e72;
        12'd0632: out <= 24'h347c7e;
        12'd0633: out <= 24'h327b8c;
        12'd0634: out <= 24'h347e9d;
        12'd0635: out <= 24'h3680ae;
        12'd0636: out <= 24'h347ebc;
        12'd0637: out <= 24'h327cc9;
        12'd0638: out <= 24'h347fda;
        12'd0639: out <= 24'h347fda;
        12'd0640: out <= 24'h378b05;
        12'd0641: out <= 24'h358a12;
        12'd0642: out <= 24'h33881f;
        12'd0643: out <= 24'h358a30;
        12'd0644: out <= 24'h378d42;
        12'd0645: out <= 24'h358c50;
        12'd0646: out <= 24'h338a5d;
        12'd0647: out <= 24'h368c6e;
        12'd0648: out <= 24'h388f80;
        12'd0649: out <= 24'h368e8d;
        12'd0650: out <= 24'h348c9a;
        12'd0651: out <= 24'h368eac;
        12'd0652: out <= 24'h3991bd;
        12'd0653: out <= 24'h378fca;
        12'd0654: out <= 24'h358dd7;
        12'd0655: out <= 24'h358dd7;
        12'd0656: out <= 24'h379a02;
        12'd0657: out <= 24'h399c14;
        12'd0658: out <= 24'h379a20;
        12'd0659: out <= 24'h36992e;
        12'd0660: out <= 24'h389c3f;
        12'd0661: out <= 24'h3a9e50;
        12'd0662: out <= 24'h389c5e;
        12'd0663: out <= 24'h369b6c;
        12'd0664: out <= 24'h389e7d;
        12'd0665: out <= 24'h3aa08e;
        12'd0666: out <= 24'h389e9b;
        12'd0667: out <= 24'h369da8;
        12'd0668: out <= 24'h39a0ba;
        12'd0669: out <= 24'h3ba2cc;
        12'd0670: out <= 24'h39a0d8;
        12'd0671: out <= 24'h39a0d8;
        12'd0672: out <= 24'h37a800;
        12'd0673: out <= 24'h39aa11;
        12'd0674: out <= 24'h3bad22;
        12'd0675: out <= 24'h3aac2f;
        12'd0676: out <= 24'h38aa3c;
        12'd0677: out <= 24'h3aac4e;
        12'd0678: out <= 24'h3caf5f;
        12'd0679: out <= 24'h3aae6c;
        12'd0680: out <= 24'h38ac7a;
        12'd0681: out <= 24'h3aae8b;
        12'd0682: out <= 24'h3db19c;
        12'd0683: out <= 24'h3bb0aa;
        12'd0684: out <= 24'h39aeb7;
        12'd0685: out <= 24'h3bb0c8;
        12'd0686: out <= 24'h3db3da;
        12'd0687: out <= 24'h3db3da;
        12'd0688: out <= 24'h3cbb00;
        12'd0689: out <= 24'h3ab90e;
        12'd0690: out <= 24'h3cbc1f;
        12'd0691: out <= 24'h3ebe30;
        12'd0692: out <= 24'h3cbc3e;
        12'd0693: out <= 24'h3abb4a;
        12'd0694: out <= 24'h3cbe5c;
        12'd0695: out <= 24'h3ec06e;
        12'd0696: out <= 24'h3cbe7b;
        12'd0697: out <= 24'h3abd88;
        12'd0698: out <= 24'h3dc099;
        12'd0699: out <= 24'h40c2aa;
        12'd0700: out <= 24'h3ec0b8;
        12'd0701: out <= 24'h3cbfc6;
        12'd0702: out <= 24'h3ec2d7;
        12'd0703: out <= 24'h3ec2d7;
        12'd0704: out <= 24'h40ce01;
        12'd0705: out <= 24'h3ecc0e;
        12'd0706: out <= 24'h3cca1c;
        12'd0707: out <= 24'h3ecc2e;
        12'd0708: out <= 24'h40cf3f;
        12'd0709: out <= 24'h3ece4c;
        12'd0710: out <= 24'h3dcc59;
        12'd0711: out <= 24'h3fce6a;
        12'd0712: out <= 24'h41d17c;
        12'd0713: out <= 24'h3fd089;
        12'd0714: out <= 24'h3dce96;
        12'd0715: out <= 24'h40d0a8;
        12'd0716: out <= 24'h42d3b9;
        12'd0717: out <= 24'h40d2c6;
        12'd0718: out <= 24'h3ed0d4;
        12'd0719: out <= 24'h3ed0d4;
        12'd0720: out <= 24'h44e002;
        12'd0721: out <= 24'h42df10;
        12'd0722: out <= 24'h40dd1d;
        12'd0723: out <= 24'h42e02e;
        12'd0724: out <= 24'h44e240;
        12'd0725: out <= 24'h42e04d;
        12'd0726: out <= 24'h41de5a;
        12'd0727: out <= 24'h44e16c;
        12'd0728: out <= 24'h46e47d;
        12'd0729: out <= 24'h44e28a;
        12'd0730: out <= 24'h42e098;
        12'd0731: out <= 24'h44e3a8;
        12'd0732: out <= 24'h46e6ba;
        12'd0733: out <= 24'h44e4c8;
        12'd0734: out <= 24'h42e2d5;
        12'd0735: out <= 24'h42e2d5;
        12'd0736: out <= 24'h48f303;
        12'd0737: out <= 24'h46f210;
        12'd0738: out <= 24'h45f01e;
        12'd0739: out <= 24'h47f230;
        12'd0740: out <= 24'h49f541;
        12'd0741: out <= 24'h47f34e;
        12'd0742: out <= 24'h45f15b;
        12'd0743: out <= 24'h48f46c;
        12'd0744: out <= 24'h4af67e;
        12'd0745: out <= 24'h48f48c;
        12'd0746: out <= 24'h46f399;
        12'd0747: out <= 24'h48f6aa;
        12'd0748: out <= 24'h4af8bb;
        12'd0749: out <= 24'h48f6c8;
        12'd0750: out <= 24'h47f5d6;
        12'd0751: out <= 24'h47f5d6;
        12'd0752: out <= 24'h48f303;
        12'd0753: out <= 24'h46f210;
        12'd0754: out <= 24'h45f01e;
        12'd0755: out <= 24'h47f230;
        12'd0756: out <= 24'h49f541;
        12'd0757: out <= 24'h47f34e;
        12'd0758: out <= 24'h45f15b;
        12'd0759: out <= 24'h48f46c;
        12'd0760: out <= 24'h4af67e;
        12'd0761: out <= 24'h48f48c;
        12'd0762: out <= 24'h46f399;
        12'd0763: out <= 24'h48f6aa;
        12'd0764: out <= 24'h4af8bb;
        12'd0765: out <= 24'h48f6c8;
        12'd0766: out <= 24'h47f5d6;
        12'd0767: out <= 24'h47f5d6;
        12'd0768: out <= 24'h2e030a;
        12'd0769: out <= 24'h2c0218;
        12'd0770: out <= 24'h2e0429;
        12'd0771: out <= 24'h30063a;
        12'd0772: out <= 24'h2f0448;
        12'd0773: out <= 24'h2d0354;
        12'd0774: out <= 24'h2f0666;
        12'd0775: out <= 24'h320878;
        12'd0776: out <= 24'h300685;
        12'd0777: out <= 24'h2e0492;
        12'd0778: out <= 24'h3006a4;
        12'd0779: out <= 24'h3209b5;
        12'd0780: out <= 24'h3008c2;
        12'd0781: out <= 24'h2e06d0;
        12'd0782: out <= 24'h3008e1;
        12'd0783: out <= 24'h3008e1;
        12'd0784: out <= 24'h2e1207;
        12'd0785: out <= 24'h301418;
        12'd0786: out <= 24'h32162a;
        12'd0787: out <= 24'h301438;
        12'd0788: out <= 24'h2f1344;
        12'd0789: out <= 24'h321656;
        12'd0790: out <= 24'h341868;
        12'd0791: out <= 24'h321674;
        12'd0792: out <= 24'h301482;
        12'd0793: out <= 24'h321794;
        12'd0794: out <= 24'h341aa5;
        12'd0795: out <= 24'h3218b2;
        12'd0796: out <= 24'h3016bf;
        12'd0797: out <= 24'h3218d0;
        12'd0798: out <= 24'h341be2;
        12'd0799: out <= 24'h341be2;
        12'd0800: out <= 24'h332408;
        12'd0801: out <= 24'h35261a;
        12'd0802: out <= 24'h332427;
        12'd0803: out <= 24'h312334;
        12'd0804: out <= 24'h332646;
        12'd0805: out <= 24'h362858;
        12'd0806: out <= 24'h342664;
        12'd0807: out <= 24'h322572;
        12'd0808: out <= 24'h342883;
        12'd0809: out <= 24'h362a94;
        12'd0810: out <= 24'h3428a2;
        12'd0811: out <= 24'h3226af;
        12'd0812: out <= 24'h3528c0;
        12'd0813: out <= 24'h372bd2;
        12'd0814: out <= 24'h352adf;
        12'd0815: out <= 24'h352adf;
        12'd0816: out <= 24'h37360a;
        12'd0817: out <= 24'h363416;
        12'd0818: out <= 24'h343324;
        12'd0819: out <= 24'h363636;
        12'd0820: out <= 24'h383847;
        12'd0821: out <= 24'h363654;
        12'd0822: out <= 24'h343562;
        12'd0823: out <= 24'h363872;
        12'd0824: out <= 24'h383a84;
        12'd0825: out <= 24'h363892;
        12'd0826: out <= 24'h34369f;
        12'd0827: out <= 24'h3639b0;
        12'd0828: out <= 24'h393cc2;
        12'd0829: out <= 24'h383ace;
        12'd0830: out <= 24'h3638dc;
        12'd0831: out <= 24'h3638dc;
        12'd0832: out <= 24'h3b480b;
        12'd0833: out <= 24'h3a4718;
        12'd0834: out <= 24'h384625;
        12'd0835: out <= 24'h3a4836;
        12'd0836: out <= 24'h3c4a48;
        12'd0837: out <= 24'h3a4956;
        12'd0838: out <= 24'h384863;
        12'd0839: out <= 24'h3a4a74;
        12'd0840: out <= 24'h3d4c85;
        12'd0841: out <= 24'h3b4b92;
        12'd0842: out <= 24'h394aa0;
        12'd0843: out <= 24'h3b4cb2;
        12'd0844: out <= 24'h394abe;
        12'd0845: out <= 24'h3848cc;
        12'd0846: out <= 24'h3a4add;
        12'd0847: out <= 24'h3a4add;
        12'd0848: out <= 24'h3c5708;
        12'd0849: out <= 24'h3e5a1a;
        12'd0850: out <= 24'h3c5826;
        12'd0851: out <= 24'h3a5634;
        12'd0852: out <= 24'h3c5945;
        12'd0853: out <= 24'h3e5c56;
        12'd0854: out <= 24'h3c5a64;
        12'd0855: out <= 24'h3a5871;
        12'd0856: out <= 24'h3d5b82;
        12'd0857: out <= 24'h405e94;
        12'd0858: out <= 24'h3e5ca1;
        12'd0859: out <= 24'h3c5aae;
        12'd0860: out <= 24'h3a58bc;
        12'd0861: out <= 24'h3c5bcd;
        12'd0862: out <= 24'h3e5ede;
        12'd0863: out <= 24'h3e5ede;
        12'd0864: out <= 24'h3c6605;
        12'd0865: out <= 24'h3e6816;
        12'd0866: out <= 24'h406a28;
        12'd0867: out <= 24'h3e6934;
        12'd0868: out <= 24'h3c6842;
        12'd0869: out <= 24'h3e6a54;
        12'd0870: out <= 24'h416c65;
        12'd0871: out <= 24'h3f6b72;
        12'd0872: out <= 24'h3d6a7f;
        12'd0873: out <= 24'h406c90;
        12'd0874: out <= 24'h426ea2;
        12'd0875: out <= 24'h406db0;
        12'd0876: out <= 24'h3e6cbd;
        12'd0877: out <= 24'h406ece;
        12'd0878: out <= 24'h4270e0;
        12'd0879: out <= 24'h4270e0;
        12'd0880: out <= 24'h407806;
        12'd0881: out <= 24'h427a18;
        12'd0882: out <= 24'h447d28;
        12'd0883: out <= 24'h427c36;
        12'd0884: out <= 24'h407a43;
        12'd0885: out <= 24'h437c54;
        12'd0886: out <= 24'h467f66;
        12'd0887: out <= 24'h447e74;
        12'd0888: out <= 24'h427c80;
        12'd0889: out <= 24'h447e92;
        12'd0890: out <= 24'h4681a3;
        12'd0891: out <= 24'h4480b0;
        12'd0892: out <= 24'h427ebe;
        12'd0893: out <= 24'h4480d0;
        12'd0894: out <= 24'h4683e0;
        12'd0895: out <= 24'h4683e0;
        12'd0896: out <= 24'h458a07;
        12'd0897: out <= 24'h478d18;
        12'd0898: out <= 24'h458c26;
        12'd0899: out <= 24'h438a32;
        12'd0900: out <= 24'h458c44;
        12'd0901: out <= 24'h488f56;
        12'd0902: out <= 24'h468e63;
        12'd0903: out <= 24'h448c70;
        12'd0904: out <= 24'h468e82;
        12'd0905: out <= 24'h489193;
        12'd0906: out <= 24'h4690a0;
        12'd0907: out <= 24'h448eae;
        12'd0908: out <= 24'h4790bf;
        12'd0909: out <= 24'h4993d0;
        12'd0910: out <= 24'h4791de;
        12'd0911: out <= 24'h4791de;
        12'd0912: out <= 24'h499e08;
        12'd0913: out <= 24'h479c16;
        12'd0914: out <= 24'h459a22;
        12'd0915: out <= 24'h489c34;
        12'd0916: out <= 24'h4a9f46;
        12'd0917: out <= 24'h489e52;
        12'd0918: out <= 24'h469c60;
        12'd0919: out <= 24'h489e72;
        12'd0920: out <= 24'h4aa183;
        12'd0921: out <= 24'h48a090;
        12'd0922: out <= 24'h469e9d;
        12'd0923: out <= 24'h48a0ae;
        12'd0924: out <= 24'h4ba3c0;
        12'd0925: out <= 24'h49a2ce;
        12'd0926: out <= 24'h47a0da;
        12'd0927: out <= 24'h47a0da;
        12'd0928: out <= 24'h49ac06;
        12'd0929: out <= 24'h47aa13;
        12'd0930: out <= 24'h49ac24;
        12'd0931: out <= 24'h4caf36;
        12'd0932: out <= 24'h4aae42;
        12'd0933: out <= 24'h48ac50;
        12'd0934: out <= 24'h4aae61;
        12'd0935: out <= 24'h4cb172;
        12'd0936: out <= 24'h4ab080;
        12'd0937: out <= 24'h48ae8d;
        12'd0938: out <= 24'h4bb09e;
        12'd0939: out <= 24'h4db3b0;
        12'd0940: out <= 24'h4bb2bd;
        12'd0941: out <= 24'h49b0ca;
        12'd0942: out <= 24'h4bb2dc;
        12'd0943: out <= 24'h4bb2dc;
        12'd0944: out <= 24'h4aba02;
        12'd0945: out <= 24'h4cbd14;
        12'd0946: out <= 24'h4ec025;
        12'd0947: out <= 24'h4cbe32;
        12'd0948: out <= 24'h4abc40;
        12'd0949: out <= 24'h4cbe50;
        12'd0950: out <= 24'h4ec162;
        12'd0951: out <= 24'h4cc070;
        12'd0952: out <= 24'h4abe7d;
        12'd0953: out <= 24'h4cc08e;
        12'd0954: out <= 24'h4fc3a0;
        12'd0955: out <= 24'h4ec2ac;
        12'd0956: out <= 24'h4cc0ba;
        12'd0957: out <= 24'h4ec2cc;
        12'd0958: out <= 24'h50c5dd;
        12'd0959: out <= 24'h50c5dd;
        12'd0960: out <= 24'h4ece03;
        12'd0961: out <= 24'h50d014;
        12'd0962: out <= 24'h4ece22;
        12'd0963: out <= 24'h4ccc30;
        12'd0964: out <= 24'h4ece41;
        12'd0965: out <= 24'h50d152;
        12'd0966: out <= 24'h4fd05f;
        12'd0967: out <= 24'h4dce6c;
        12'd0968: out <= 24'h4fd07e;
        12'd0969: out <= 24'h51d390;
        12'd0970: out <= 24'h4fd29c;
        12'd0971: out <= 24'h4ed0aa;
        12'd0972: out <= 24'h50d2bb;
        12'd0973: out <= 24'h52d5cc;
        12'd0974: out <= 24'h50d4da;
        12'd0975: out <= 24'h50d4da;
        12'd0976: out <= 24'h52e004;
        12'd0977: out <= 24'h50de12;
        12'd0978: out <= 24'h4edc1f;
        12'd0979: out <= 24'h50de30;
        12'd0980: out <= 24'h52e142;
        12'd0981: out <= 24'h50e04f;
        12'd0982: out <= 24'h4fde5c;
        12'd0983: out <= 24'h52e06e;
        12'd0984: out <= 24'h54e37f;
        12'd0985: out <= 24'h52e28c;
        12'd0986: out <= 24'h50e09a;
        12'd0987: out <= 24'h52e2ab;
        12'd0988: out <= 24'h54e5bc;
        12'd0989: out <= 24'h52e4ca;
        12'd0990: out <= 24'h50e2d7;
        12'd0991: out <= 24'h50e2d7;
        12'd0992: out <= 24'h56f206;
        12'd0993: out <= 24'h54f012;
        12'd0994: out <= 24'h53ef20;
        12'd0995: out <= 24'h55f232;
        12'd0996: out <= 24'h57f443;
        12'd0997: out <= 24'h55f250;
        12'd0998: out <= 24'h53f05d;
        12'd0999: out <= 24'h56f36e;
        12'd1000: out <= 24'h58f680;
        12'd1001: out <= 24'h56f48e;
        12'd1002: out <= 24'h54f29b;
        12'd1003: out <= 24'h56f5ac;
        12'd1004: out <= 24'h58f8be;
        12'd1005: out <= 24'h56f6ca;
        12'd1006: out <= 24'h55f4d8;
        12'd1007: out <= 24'h55f4d8;
        12'd1008: out <= 24'h56f206;
        12'd1009: out <= 24'h54f012;
        12'd1010: out <= 24'h53ef20;
        12'd1011: out <= 24'h55f232;
        12'd1012: out <= 24'h57f443;
        12'd1013: out <= 24'h55f250;
        12'd1014: out <= 24'h53f05d;
        12'd1015: out <= 24'h56f36e;
        12'd1016: out <= 24'h58f680;
        12'd1017: out <= 24'h56f48e;
        12'd1018: out <= 24'h54f29b;
        12'd1019: out <= 24'h56f5ac;
        12'd1020: out <= 24'h58f8be;
        12'd1021: out <= 24'h56f6ca;
        12'd1022: out <= 24'h55f4d8;
        12'd1023: out <= 24'h55f4d8;
        12'd1024: out <= 24'h400610;
        12'd1025: out <= 24'h3e041e;
        12'd1026: out <= 24'h3c032b;
        12'd1027: out <= 24'h3e063c;
        12'd1028: out <= 24'h41084e;
        12'd1029: out <= 24'h3f065b;
        12'd1030: out <= 24'h3d0568;
        12'd1031: out <= 24'h40087a;
        12'd1032: out <= 24'h420a8b;
        12'd1033: out <= 24'h400898;
        12'd1034: out <= 24'h3e06a6;
        12'd1035: out <= 24'h4008b7;
        12'd1036: out <= 24'h420bc8;
        12'd1037: out <= 24'h400ad6;
        12'd1038: out <= 24'h3e08e3;
        12'd1039: out <= 24'h3e08e3;
        12'd1040: out <= 24'h40140d;
        12'd1041: out <= 24'h42171e;
        12'd1042: out <= 24'h40162c;
        12'd1043: out <= 24'h3e143a;
        12'd1044: out <= 24'h41164b;
        12'd1045: out <= 24'h44195c;
        12'd1046: out <= 24'h42186a;
        12'd1047: out <= 24'h401676;
        12'd1048: out <= 24'h421888;
        12'd1049: out <= 24'h441b9a;
        12'd1050: out <= 24'h4219a7;
        12'd1051: out <= 24'h4017b4;
        12'd1052: out <= 24'h421ac5;
        12'd1053: out <= 24'h441cd6;
        12'd1054: out <= 24'h421ae4;
        12'd1055: out <= 24'h421ae4;
        12'd1056: out <= 24'h41230a;
        12'd1057: out <= 24'h43261c;
        12'd1058: out <= 24'h45282d;
        12'd1059: out <= 24'h43263a;
        12'd1060: out <= 24'h412548;
        12'd1061: out <= 24'h44285a;
        12'd1062: out <= 24'h462a6b;
        12'd1063: out <= 24'h442878;
        12'd1064: out <= 24'h422785;
        12'd1065: out <= 24'h442a96;
        12'd1066: out <= 24'h462ca8;
        12'd1067: out <= 24'h442ab5;
        12'd1068: out <= 24'h4328c2;
        12'd1069: out <= 24'h452ad4;
        12'd1070: out <= 24'h472de5;
        12'd1071: out <= 24'h472de5;
        12'd1072: out <= 24'h45360c;
        12'd1073: out <= 24'h443418;
        12'd1074: out <= 24'h46362a;
        12'd1075: out <= 24'h48393c;
        12'd1076: out <= 24'h463849;
        12'd1077: out <= 24'h443656;
        12'd1078: out <= 24'h463868;
        12'd1079: out <= 24'h483b79;
        12'd1080: out <= 24'h463a86;
        12'd1081: out <= 24'h443894;
        12'd1082: out <= 24'h463aa5;
        12'd1083: out <= 24'h483db6;
        12'd1084: out <= 24'h473bc4;
        12'd1085: out <= 24'h4639d0;
        12'd1086: out <= 24'h483ce2;
        12'd1087: out <= 24'h483ce2;
        12'd1088: out <= 24'h49480d;
        12'd1089: out <= 24'h48461a;
        12'd1090: out <= 24'h464527;
        12'd1091: out <= 24'h484838;
        12'd1092: out <= 24'h4a4a4a;
        12'd1093: out <= 24'h484858;
        12'd1094: out <= 24'h464765;
        12'd1095: out <= 24'h484a76;
        12'd1096: out <= 24'h4b4c87;
        12'd1097: out <= 24'h494a94;
        12'd1098: out <= 24'h4749a2;
        12'd1099: out <= 24'h494cb4;
        12'd1100: out <= 24'h4b4ec5;
        12'd1101: out <= 24'h4a4cd2;
        12'd1102: out <= 24'h484adf;
        12'd1103: out <= 24'h484adf;
        12'd1104: out <= 24'h4a560a;
        12'd1105: out <= 24'h4c591c;
        12'd1106: out <= 24'h4a5828;
        12'd1107: out <= 24'h485636;
        12'd1108: out <= 24'h4a5847;
        12'd1109: out <= 24'h4c5b58;
        12'd1110: out <= 24'h4a5a66;
        12'd1111: out <= 24'h485873;
        12'd1112: out <= 24'h4b5a84;
        12'd1113: out <= 24'h4e5d96;
        12'd1114: out <= 24'h4c5ca3;
        12'd1115: out <= 24'h4a5ab0;
        12'd1116: out <= 24'h4c5cc2;
        12'd1117: out <= 24'h4e5fd4;
        12'd1118: out <= 24'h4c5de0;
        12'd1119: out <= 24'h4c5de0;
        12'd1120: out <= 24'h4a6507;
        12'd1121: out <= 24'h4c6818;
        12'd1122: out <= 24'h4e6a2a;
        12'd1123: out <= 24'h4c6837;
        12'd1124: out <= 24'h4a6744;
        12'd1125: out <= 24'h4c6a56;
        12'd1126: out <= 24'h4f6c67;
        12'd1127: out <= 24'h4d6a74;
        12'd1128: out <= 24'h4b6981;
        12'd1129: out <= 24'h4e6c92;
        12'd1130: out <= 24'h506ea4;
        12'd1131: out <= 24'h4e6cb2;
        12'd1132: out <= 24'h4c6bbf;
        12'd1133: out <= 24'h4e6ed0;
        12'd1134: out <= 24'h5070e2;
        12'd1135: out <= 24'h5070e2;
        12'd1136: out <= 24'h4e7808;
        12'd1137: out <= 24'h507a1a;
        12'd1138: out <= 24'h527c2b;
        12'd1139: out <= 24'h507b38;
        12'd1140: out <= 24'h4e7a45;
        12'd1141: out <= 24'h517c56;
        12'd1142: out <= 24'h547e68;
        12'd1143: out <= 24'h527d76;
        12'd1144: out <= 24'h507c82;
        12'd1145: out <= 24'h527e94;
        12'd1146: out <= 24'h5480a5;
        12'd1147: out <= 24'h527fb2;
        12'd1148: out <= 24'h507ec0;
        12'd1149: out <= 24'h5280d2;
        12'd1150: out <= 24'h5482e3;
        12'd1151: out <= 24'h5482e3;
        12'd1152: out <= 24'h538a09;
        12'd1153: out <= 24'h558c1a;
        12'd1154: out <= 24'h578f2c;
        12'd1155: out <= 24'h558e39;
        12'd1156: out <= 24'h538c46;
        12'd1157: out <= 24'h568e58;
        12'd1158: out <= 24'h589169;
        12'd1159: out <= 24'h569076;
        12'd1160: out <= 24'h548e84;
        12'd1161: out <= 24'h569095;
        12'd1162: out <= 24'h5893a6;
        12'd1163: out <= 24'h5692b4;
        12'd1164: out <= 24'h5590c1;
        12'd1165: out <= 24'h5792d2;
        12'd1166: out <= 24'h5995e4;
        12'd1167: out <= 24'h5995e4;
        12'd1168: out <= 24'h579d0a;
        12'd1169: out <= 24'h559b18;
        12'd1170: out <= 24'h579e29;
        12'd1171: out <= 24'h5aa03a;
        12'd1172: out <= 24'h589e48;
        12'd1173: out <= 24'h569d54;
        12'd1174: out <= 24'h58a066;
        12'd1175: out <= 24'h5aa278;
        12'd1176: out <= 24'h58a085;
        12'd1177: out <= 24'h569f92;
        12'd1178: out <= 24'h58a2a3;
        12'd1179: out <= 24'h5aa4b4;
        12'd1180: out <= 24'h59a2c2;
        12'd1181: out <= 24'h57a1d0;
        12'd1182: out <= 24'h59a4e1;
        12'd1183: out <= 24'h59a4e1;
        12'd1184: out <= 24'h5bb00b;
        12'd1185: out <= 24'h59ae18;
        12'd1186: out <= 24'h57ac26;
        12'd1187: out <= 24'h5aae38;
        12'd1188: out <= 24'h5cb149;
        12'd1189: out <= 24'h5ab056;
        12'd1190: out <= 24'h58ae63;
        12'd1191: out <= 24'h5ab074;
        12'd1192: out <= 24'h5db386;
        12'd1193: out <= 24'h5bb293;
        12'd1194: out <= 24'h59b0a0;
        12'd1195: out <= 24'h5bb2b2;
        12'd1196: out <= 24'h5db5c3;
        12'd1197: out <= 24'h5bb4d0;
        12'd1198: out <= 24'h59b2de;
        12'd1199: out <= 24'h59b2de;
        12'd1200: out <= 24'h5cbe08;
        12'd1201: out <= 24'h5ec11a;
        12'd1202: out <= 24'h5cbf27;
        12'd1203: out <= 24'h5abd34;
        12'd1204: out <= 24'h5cc046;
        12'd1205: out <= 24'h5ec257;
        12'd1206: out <= 24'h5cc064;
        12'd1207: out <= 24'h5abf72;
        12'd1208: out <= 24'h5dc283;
        12'd1209: out <= 24'h5fc494;
        12'd1210: out <= 24'h5dc2a2;
        12'd1211: out <= 24'h5cc1ae;
        12'd1212: out <= 24'h5ec4c0;
        12'd1213: out <= 24'h60c6d2;
        12'd1214: out <= 24'h5ec4df;
        12'd1215: out <= 24'h5ec4df;
        12'd1216: out <= 24'h5ccd05;
        12'd1217: out <= 24'h5ed016;
        12'd1218: out <= 24'h60d228;
        12'd1219: out <= 24'h5ed036;
        12'd1220: out <= 24'h5cce43;
        12'd1221: out <= 24'h5ed054;
        12'd1222: out <= 24'h61d365;
        12'd1223: out <= 24'h5fd272;
        12'd1224: out <= 24'h5dd080;
        12'd1225: out <= 24'h5fd292;
        12'd1226: out <= 24'h61d5a3;
        12'd1227: out <= 24'h60d4b0;
        12'd1228: out <= 24'h5ed2bd;
        12'd1229: out <= 24'h60d4ce;
        12'd1230: out <= 24'h62d7e0;
        12'd1231: out <= 24'h62d7e0;
        12'd1232: out <= 24'h60e006;
        12'd1233: out <= 24'h5ede14;
        12'd1234: out <= 24'h60e025;
        12'd1235: out <= 24'h62e236;
        12'd1236: out <= 24'h60e044;
        12'd1237: out <= 24'h5edf51;
        12'd1238: out <= 24'h61e262;
        12'd1239: out <= 24'h64e474;
        12'd1240: out <= 24'h62e281;
        12'd1241: out <= 24'h60e18e;
        12'd1242: out <= 24'h62e4a0;
        12'd1243: out <= 24'h64e6b2;
        12'd1244: out <= 24'h62e4be;
        12'd1245: out <= 24'h60e3cc;
        12'd1246: out <= 24'h62e6dd;
        12'd1247: out <= 24'h62e6dd;
        12'd1248: out <= 24'h64f208;
        12'd1249: out <= 24'h62f015;
        12'd1250: out <= 24'h61ee22;
        12'd1251: out <= 24'h63f034;
        12'd1252: out <= 24'h65f345;
        12'd1253: out <= 24'h63f252;
        12'd1254: out <= 24'h61f05f;
        12'd1255: out <= 24'h64f270;
        12'd1256: out <= 24'h66f582;
        12'd1257: out <= 24'h64f490;
        12'd1258: out <= 24'h62f29d;
        12'd1259: out <= 24'h64f4ae;
        12'd1260: out <= 24'h66f7c0;
        12'd1261: out <= 24'h64f6cd;
        12'd1262: out <= 24'h63f4da;
        12'd1263: out <= 24'h63f4da;
        12'd1264: out <= 24'h64f208;
        12'd1265: out <= 24'h62f015;
        12'd1266: out <= 24'h61ee22;
        12'd1267: out <= 24'h63f034;
        12'd1268: out <= 24'h65f345;
        12'd1269: out <= 24'h63f252;
        12'd1270: out <= 24'h61f05f;
        12'd1271: out <= 24'h64f270;
        12'd1272: out <= 24'h66f582;
        12'd1273: out <= 24'h64f490;
        12'd1274: out <= 24'h62f29d;
        12'd1275: out <= 24'h64f4ae;
        12'd1276: out <= 24'h66f7c0;
        12'd1277: out <= 24'h64f6cd;
        12'd1278: out <= 24'h63f4da;
        12'd1279: out <= 24'h63f4da;
        12'd1280: out <= 24'h4e0612;
        12'd1281: out <= 24'h4c0420;
        12'd1282: out <= 24'h4a022d;
        12'd1283: out <= 24'h4c053e;
        12'd1284: out <= 24'h4f0850;
        12'd1285: out <= 24'h4d065d;
        12'd1286: out <= 24'h4b046a;
        12'd1287: out <= 24'h4e077c;
        12'd1288: out <= 24'h500a8d;
        12'd1289: out <= 24'h4e089a;
        12'd1290: out <= 24'h4c06a8;
        12'd1291: out <= 24'h4e08ba;
        12'd1292: out <= 24'h500aca;
        12'd1293: out <= 24'h4e09d8;
        12'd1294: out <= 24'h4c08e5;
        12'd1295: out <= 24'h4c08e5;
        12'd1296: out <= 24'h521814;
        12'd1297: out <= 24'h501620;
        12'd1298: out <= 24'h4e152e;
        12'd1299: out <= 24'h511840;
        12'd1300: out <= 24'h541a51;
        12'd1301: out <= 24'h52185e;
        12'd1302: out <= 24'h50176c;
        12'd1303: out <= 24'h521a7c;
        12'd1304: out <= 24'h541c8e;
        12'd1305: out <= 24'h521a9c;
        12'd1306: out <= 24'h5018a9;
        12'd1307: out <= 24'h521bba;
        12'd1308: out <= 24'h541ecc;
        12'd1309: out <= 24'h521cd8;
        12'd1310: out <= 24'h501ae6;
        12'd1311: out <= 24'h501ae6;
        12'd1312: out <= 24'h532610;
        12'd1313: out <= 24'h51251e;
        12'd1314: out <= 24'h53282f;
        12'd1315: out <= 24'h562a40;
        12'd1316: out <= 24'h54284e;
        12'd1317: out <= 24'h52275c;
        12'd1318: out <= 24'h542a6d;
        12'd1319: out <= 24'h562c7e;
        12'd1320: out <= 24'h542a8b;
        12'd1321: out <= 24'h522998;
        12'd1322: out <= 24'h542caa;
        12'd1323: out <= 24'h562ebc;
        12'd1324: out <= 24'h552cc8;
        12'd1325: out <= 24'h532ad6;
        12'd1326: out <= 24'h552ce7;
        12'd1327: out <= 24'h552ce7;
        12'd1328: out <= 24'h53350e;
        12'd1329: out <= 24'h56381f;
        12'd1330: out <= 24'h583a30;
        12'd1331: out <= 24'h56383e;
        12'd1332: out <= 24'h54374b;
        12'd1333: out <= 24'h563a5c;
        12'd1334: out <= 24'h583c6e;
        12'd1335: out <= 24'h563a7b;
        12'd1336: out <= 24'h543988;
        12'd1337: out <= 24'h563c9a;
        12'd1338: out <= 24'h583eab;
        12'd1339: out <= 24'h563cb8;
        12'd1340: out <= 24'h553ac6;
        12'd1341: out <= 24'h583dd7;
        12'd1342: out <= 24'h5a40e8;
        12'd1343: out <= 24'h5a40e8;
        12'd1344: out <= 24'h57480f;
        12'd1345: out <= 24'h5a4a20;
        12'd1346: out <= 24'h58482e;
        12'd1347: out <= 24'h56473a;
        12'd1348: out <= 24'h584a4c;
        12'd1349: out <= 24'h5a4c5e;
        12'd1350: out <= 24'h584a6b;
        12'd1351: out <= 24'h564978;
        12'd1352: out <= 24'h594c89;
        12'd1353: out <= 24'h5b4e9a;
        12'd1354: out <= 24'h594ca8;
        12'd1355: out <= 24'h574bb6;
        12'd1356: out <= 24'h594ec7;
        12'd1357: out <= 24'h5c50d8;
        12'd1358: out <= 24'h5a4ee6;
        12'd1359: out <= 24'h5a4ee6;
        12'd1360: out <= 24'h5c5a10;
        12'd1361: out <= 24'h5a581e;
        12'd1362: out <= 24'h58572a;
        12'd1363: out <= 24'h5a5a3c;
        12'd1364: out <= 24'h5c5c4d;
        12'd1365: out <= 24'h5a5a5a;
        12'd1366: out <= 24'h585968;
        12'd1367: out <= 24'h5a5c7a;
        12'd1368: out <= 24'h5d5e8a;
        12'd1369: out <= 24'h5c5c98;
        12'd1370: out <= 24'h5a5ba5;
        12'd1371: out <= 24'h5c5eb6;
        12'd1372: out <= 24'h5e60c8;
        12'd1373: out <= 24'h5c5ed6;
        12'd1374: out <= 24'h5a5ce2;
        12'd1375: out <= 24'h5a5ce2;
        12'd1376: out <= 24'h5c680d;
        12'd1377: out <= 24'h5a671a;
        12'd1378: out <= 24'h5c6a2c;
        12'd1379: out <= 24'h5e6c3d;
        12'd1380: out <= 24'h5c6a4a;
        12'd1381: out <= 24'h5a6958;
        12'd1382: out <= 24'h5d6c69;
        12'd1383: out <= 24'h5f6e7a;
        12'd1384: out <= 24'h5d6c88;
        12'd1385: out <= 24'h5c6b94;
        12'd1386: out <= 24'h5e6ea6;
        12'd1387: out <= 24'h6070b8;
        12'd1388: out <= 24'h5e6ec5;
        12'd1389: out <= 24'h5c6cd2;
        12'd1390: out <= 24'h5e6fe4;
        12'd1391: out <= 24'h5e6fe4;
        12'd1392: out <= 24'h5c770a;
        12'd1393: out <= 24'h5e7a1c;
        12'd1394: out <= 24'h607c2d;
        12'd1395: out <= 24'h5e7a3a;
        12'd1396: out <= 24'h5c7947;
        12'd1397: out <= 24'h5f7c58;
        12'd1398: out <= 24'h627e6a;
        12'd1399: out <= 24'h607c78;
        12'd1400: out <= 24'h5e7b84;
        12'd1401: out <= 24'h607e96;
        12'd1402: out <= 24'h6280a8;
        12'd1403: out <= 24'h607eb4;
        12'd1404: out <= 24'h5e7dc2;
        12'd1405: out <= 24'h6080d4;
        12'd1406: out <= 24'h6282e5;
        12'd1407: out <= 24'h6282e5;
        12'd1408: out <= 24'h618a0b;
        12'd1409: out <= 24'h638c1c;
        12'd1410: out <= 24'h658e2e;
        12'd1411: out <= 24'h638d3b;
        12'd1412: out <= 24'h618c48;
        12'd1413: out <= 24'h648e5a;
        12'd1414: out <= 24'h66906b;
        12'd1415: out <= 24'h648f78;
        12'd1416: out <= 24'h628e86;
        12'd1417: out <= 24'h649098;
        12'd1418: out <= 24'h6692a8;
        12'd1419: out <= 24'h6491b6;
        12'd1420: out <= 24'h6390c3;
        12'd1421: out <= 24'h6592d4;
        12'd1422: out <= 24'h6794e6;
        12'd1423: out <= 24'h6794e6;
        12'd1424: out <= 24'h659c0c;
        12'd1425: out <= 24'h689f1e;
        12'd1426: out <= 24'h6aa22f;
        12'd1427: out <= 24'h68a03c;
        12'd1428: out <= 24'h669e4a;
        12'd1429: out <= 24'h68a05a;
        12'd1430: out <= 24'h6aa36c;
        12'd1431: out <= 24'h68a27a;
        12'd1432: out <= 24'h66a087;
        12'd1433: out <= 24'h649e94;
        12'd1434: out <= 24'h66a1a6;
        12'd1435: out <= 24'h68a4b6;
        12'd1436: out <= 24'h67a2c4;
        12'd1437: out <= 24'h65a0d2;
        12'd1438: out <= 24'h67a3e3;
        12'd1439: out <= 24'h67a3e3;
        12'd1440: out <= 24'h69b00d;
        12'd1441: out <= 24'h6cb21e;
        12'd1442: out <= 24'h6ab02c;
        12'd1443: out <= 24'h68ae3a;
        12'd1444: out <= 24'h6ab04b;
        12'd1445: out <= 24'h6cb35c;
        12'd1446: out <= 24'h6ab269;
        12'd1447: out <= 24'h68b076;
        12'd1448: out <= 24'h6bb288;
        12'd1449: out <= 24'h69b196;
        12'd1450: out <= 24'h67b0a2;
        12'd1451: out <= 24'h69b2b4;
        12'd1452: out <= 24'h6bb4c5;
        12'd1453: out <= 24'h69b3d2;
        12'd1454: out <= 24'h67b2e0;
        12'd1455: out <= 24'h67b2e0;
        12'd1456: out <= 24'h6ec20e;
        12'd1457: out <= 24'h6cc01c;
        12'd1458: out <= 24'h6abe29;
        12'd1459: out <= 24'h6cc03a;
        12'd1460: out <= 24'h6ec34c;
        12'd1461: out <= 24'h6cc259;
        12'd1462: out <= 24'h6ac066;
        12'd1463: out <= 24'h6cc278;
        12'd1464: out <= 24'h6fc589;
        12'd1465: out <= 24'h6dc496;
        12'd1466: out <= 24'h6bc2a4;
        12'd1467: out <= 24'h6ec4b5;
        12'd1468: out <= 24'h70c7c6;
        12'd1469: out <= 24'h6ec6d4;
        12'd1470: out <= 24'h6cc4e1;
        12'd1471: out <= 24'h6cc4e1;
        12'd1472: out <= 24'h6ed00c;
        12'd1473: out <= 24'h6cce18;
        12'd1474: out <= 24'h6ed12a;
        12'd1475: out <= 24'h70d43c;
        12'd1476: out <= 24'h6ed249;
        12'd1477: out <= 24'h6cd056;
        12'd1478: out <= 24'h6fd267;
        12'd1479: out <= 24'h71d578;
        12'd1480: out <= 24'h6fd486;
        12'd1481: out <= 24'h6dd294;
        12'd1482: out <= 24'h6fd4a5;
        12'd1483: out <= 24'h72d7b6;
        12'd1484: out <= 24'h70d6c4;
        12'd1485: out <= 24'h6ed4d0;
        12'd1486: out <= 24'h70d6e2;
        12'd1487: out <= 24'h70d6e2;
        12'd1488: out <= 24'h6edf08;
        12'd1489: out <= 24'h70e21a;
        12'd1490: out <= 24'h72e42b;
        12'd1491: out <= 24'h70e238;
        12'd1492: out <= 24'h6ee046;
        12'd1493: out <= 24'h70e258;
        12'd1494: out <= 24'h73e568;
        12'd1495: out <= 24'h72e476;
        12'd1496: out <= 24'h70e283;
        12'd1497: out <= 24'h72e494;
        12'd1498: out <= 24'h74e7a6;
        12'd1499: out <= 24'h72e6b4;
        12'd1500: out <= 24'h70e4c0;
        12'd1501: out <= 24'h72e6d2;
        12'd1502: out <= 24'h74e9e3;
        12'd1503: out <= 24'h74e9e3;
        12'd1504: out <= 24'h72f20a;
        12'd1505: out <= 24'h74f41b;
        12'd1506: out <= 24'h73f228;
        12'd1507: out <= 24'h71f036;
        12'd1508: out <= 24'h73f247;
        12'd1509: out <= 24'h75f558;
        12'd1510: out <= 24'h73f466;
        12'd1511: out <= 24'h72f272;
        12'd1512: out <= 24'h74f484;
        12'd1513: out <= 24'h76f796;
        12'd1514: out <= 24'h74f6a3;
        12'd1515: out <= 24'h72f4b0;
        12'd1516: out <= 24'h74f6c2;
        12'd1517: out <= 24'h76f9d3;
        12'd1518: out <= 24'h75f8e0;
        12'd1519: out <= 24'h75f8e0;
        12'd1520: out <= 24'h72f20a;
        12'd1521: out <= 24'h74f41b;
        12'd1522: out <= 24'h73f228;
        12'd1523: out <= 24'h71f036;
        12'd1524: out <= 24'h73f247;
        12'd1525: out <= 24'h75f558;
        12'd1526: out <= 24'h73f466;
        12'd1527: out <= 24'h72f272;
        12'd1528: out <= 24'h74f484;
        12'd1529: out <= 24'h76f796;
        12'd1530: out <= 24'h74f6a3;
        12'd1531: out <= 24'h72f4b0;
        12'd1532: out <= 24'h74f6c2;
        12'd1533: out <= 24'h76f9d3;
        12'd1534: out <= 24'h75f8e0;
        12'd1535: out <= 24'h75f8e0;
        12'd1536: out <= 24'h5c0514;
        12'd1537: out <= 24'h5a0422;
        12'd1538: out <= 24'h58022f;
        12'd1539: out <= 24'h5a0440;
        12'd1540: out <= 24'h5d0752;
        12'd1541: out <= 24'h5b065f;
        12'd1542: out <= 24'h59046c;
        12'd1543: out <= 24'h5c067e;
        12'd1544: out <= 24'h5e098f;
        12'd1545: out <= 24'h5c079c;
        12'd1546: out <= 24'h5a05aa;
        12'd1547: out <= 24'h5c08bc;
        12'd1548: out <= 24'h5e0acd;
        12'd1549: out <= 24'h5c08da;
        12'd1550: out <= 24'h5a07e7;
        12'd1551: out <= 24'h5a07e7;
        12'd1552: out <= 24'h601816;
        12'd1553: out <= 24'h5e1622;
        12'd1554: out <= 24'h5c1430;
        12'd1555: out <= 24'h5f1742;
        12'd1556: out <= 24'h621a53;
        12'd1557: out <= 24'h601860;
        12'd1558: out <= 24'h5e166e;
        12'd1559: out <= 24'h60197e;
        12'd1560: out <= 24'h621c90;
        12'd1561: out <= 24'h601a9e;
        12'd1562: out <= 24'h5e18ab;
        12'd1563: out <= 24'h601abc;
        12'd1564: out <= 24'h621dce;
        12'd1565: out <= 24'h601bdb;
        12'd1566: out <= 24'h5e1ae8;
        12'd1567: out <= 24'h5e1ae8;
        12'd1568: out <= 24'h652a17;
        12'd1569: out <= 24'h632824;
        12'd1570: out <= 24'h612731;
        12'd1571: out <= 24'h642a42;
        12'd1572: out <= 24'h662c54;
        12'd1573: out <= 24'h642a62;
        12'd1574: out <= 24'h62296f;
        12'd1575: out <= 24'h642c80;
        12'd1576: out <= 24'h662e91;
        12'd1577: out <= 24'h642c9e;
        12'd1578: out <= 24'h622bac;
        12'd1579: out <= 24'h642ebe;
        12'd1580: out <= 24'h6730cf;
        12'd1581: out <= 24'h652edc;
        12'd1582: out <= 24'h632ce9;
        12'd1583: out <= 24'h632ce9;
        12'd1584: out <= 24'h653814;
        12'd1585: out <= 24'h683b26;
        12'd1586: out <= 24'h663a32;
        12'd1587: out <= 24'h643840;
        12'd1588: out <= 24'h663a51;
        12'd1589: out <= 24'h683d62;
        12'd1590: out <= 24'h663c70;
        12'd1591: out <= 24'h643a7d;
        12'd1592: out <= 24'h663c8e;
        12'd1593: out <= 24'h683fa0;
        12'd1594: out <= 24'h663ead;
        12'd1595: out <= 24'h643cba;
        12'd1596: out <= 24'h673ecc;
        12'd1597: out <= 24'h6a41de;
        12'd1598: out <= 24'h683fea;
        12'd1599: out <= 24'h683fea;
        12'd1600: out <= 24'h654711;
        12'd1601: out <= 24'h684a22;
        12'd1602: out <= 24'h6a4c34;
        12'd1603: out <= 24'h684a41;
        12'd1604: out <= 24'h66494e;
        12'd1605: out <= 24'h684c60;
        12'd1606: out <= 24'h6a4e71;
        12'd1607: out <= 24'h684c7e;
        12'd1608: out <= 24'h674b8b;
        12'd1609: out <= 24'h694e9c;
        12'd1610: out <= 24'h6b50ae;
        12'd1611: out <= 24'h694ebc;
        12'd1612: out <= 24'h674dc9;
        12'd1613: out <= 24'h6a50da;
        12'd1614: out <= 24'h6c52ec;
        12'd1615: out <= 24'h6c52ec;
        12'd1616: out <= 24'h6a5a12;
        12'd1617: out <= 24'h685820;
        12'd1618: out <= 24'h6a5a31;
        12'd1619: out <= 24'h6c5d42;
        12'd1620: out <= 24'h6a5c4f;
        12'd1621: out <= 24'h685a5c;
        12'd1622: out <= 24'h6a5c6e;
        12'd1623: out <= 24'h6c5f80;
        12'd1624: out <= 24'h6b5e8c;
        12'd1625: out <= 24'h6a5c9a;
        12'd1626: out <= 24'h6c5eab;
        12'd1627: out <= 24'h6e61bc;
        12'd1628: out <= 24'h6c60ca;
        12'd1629: out <= 24'h6a5ed8;
        12'd1630: out <= 24'h6c60e9;
        12'd1631: out <= 24'h6c60e9;
        12'd1632: out <= 24'h6e6c13;
        12'd1633: out <= 24'h6c6a20;
        12'd1634: out <= 24'h6a692e;
        12'd1635: out <= 24'h6c6c3f;
        12'd1636: out <= 24'h6f6e50;
        12'd1637: out <= 24'h6d6c5e;
        12'd1638: out <= 24'h6b6b6b;
        12'd1639: out <= 24'h6d6e7c;
        12'd1640: out <= 24'h6f708e;
        12'd1641: out <= 24'h6e6e9b;
        12'd1642: out <= 24'h6c6da8;
        12'd1643: out <= 24'h6e70ba;
        12'd1644: out <= 24'h7072cb;
        12'd1645: out <= 24'h6e70d8;
        12'd1646: out <= 24'h6c6ee6;
        12'd1647: out <= 24'h6c6ee6;
        12'd1648: out <= 24'h6e7a10;
        12'd1649: out <= 24'h707d22;
        12'd1650: out <= 24'h6e7c2f;
        12'd1651: out <= 24'h6c7a3c;
        12'd1652: out <= 24'h6f7c4d;
        12'd1653: out <= 24'h727f5e;
        12'd1654: out <= 24'h707e6c;
        12'd1655: out <= 24'h6e7c7a;
        12'd1656: out <= 24'h707e8b;
        12'd1657: out <= 24'h72819c;
        12'd1658: out <= 24'h7080aa;
        12'd1659: out <= 24'h6e7eb6;
        12'd1660: out <= 24'h7080c8;
        12'd1661: out <= 24'h7283da;
        12'd1662: out <= 24'h7081e7;
        12'd1663: out <= 24'h7081e7;
        12'd1664: out <= 24'h6f890d;
        12'd1665: out <= 24'h718c1e;
        12'd1666: out <= 24'h738e30;
        12'd1667: out <= 24'h718c3d;
        12'd1668: out <= 24'h6f8b4a;
        12'd1669: out <= 24'h728e5c;
        12'd1670: out <= 24'h74906d;
        12'd1671: out <= 24'h728e7a;
        12'd1672: out <= 24'h708d88;
        12'd1673: out <= 24'h72909a;
        12'd1674: out <= 24'h7492ab;
        12'd1675: out <= 24'h7290b8;
        12'd1676: out <= 24'h718fc5;
        12'd1677: out <= 24'h7392d6;
        12'd1678: out <= 24'h7594e8;
        12'd1679: out <= 24'h7594e8;
        12'd1680: out <= 24'h739c0e;
        12'd1681: out <= 24'h769e20;
        12'd1682: out <= 24'h78a131;
        12'd1683: out <= 24'h769f3e;
        12'd1684: out <= 24'h749e4c;
        12'd1685: out <= 24'h76a05c;
        12'd1686: out <= 24'h78a26e;
        12'd1687: out <= 24'h76a17c;
        12'd1688: out <= 24'h74a089;
        12'd1689: out <= 24'h729e96;
        12'd1690: out <= 24'h74a0a8;
        12'd1691: out <= 24'h76a3b9;
        12'd1692: out <= 24'h75a2c6;
        12'd1693: out <= 24'h73a0d4;
        12'd1694: out <= 24'h75a2e5;
        12'd1695: out <= 24'h75a2e5;
        12'd1696: out <= 24'h77af0f;
        12'd1697: out <= 24'h7ab220;
        12'd1698: out <= 24'h7cb432;
        12'd1699: out <= 24'h7ab240;
        12'd1700: out <= 24'h78b04d;
        12'd1701: out <= 24'h7ab25e;
        12'd1702: out <= 24'h7cb56f;
        12'd1703: out <= 24'h7ab47c;
        12'd1704: out <= 24'h79b28a;
        12'd1705: out <= 24'h77b098;
        12'd1706: out <= 24'h75afa5;
        12'd1707: out <= 24'h77b2b6;
        12'd1708: out <= 24'h79b4c7;
        12'd1709: out <= 24'h77b2d4;
        12'd1710: out <= 24'h75b1e2;
        12'd1711: out <= 24'h75b1e2;
        12'd1712: out <= 24'h7cc210;
        12'd1713: out <= 24'h7ac01e;
        12'd1714: out <= 24'h7cc22f;
        12'd1715: out <= 24'h7ec440;
        12'd1716: out <= 24'h7cc24e;
        12'd1717: out <= 24'h7ac15b;
        12'd1718: out <= 24'h7cc46c;
        12'd1719: out <= 24'h7ec67e;
        12'd1720: out <= 24'h7dc48b;
        12'd1721: out <= 24'h7bc398;
        12'd1722: out <= 24'h79c2a6;
        12'd1723: out <= 24'h7cc4b8;
        12'd1724: out <= 24'h7ec6c8;
        12'd1725: out <= 24'h7cc5d6;
        12'd1726: out <= 24'h7ac4e3;
        12'd1727: out <= 24'h7ac4e3;
        12'd1728: out <= 24'h80d412;
        12'd1729: out <= 24'h7ed21f;
        12'd1730: out <= 24'h7cd02c;
        12'd1731: out <= 24'h7ed23e;
        12'd1732: out <= 24'h81d54f;
        12'd1733: out <= 24'h7fd45c;
        12'd1734: out <= 24'h7dd269;
        12'd1735: out <= 24'h7fd47a;
        12'd1736: out <= 24'h81d78c;
        12'd1737: out <= 24'h7fd69a;
        12'd1738: out <= 24'h7dd4a7;
        12'd1739: out <= 24'h80d6b8;
        12'd1740: out <= 24'h82d9ca;
        12'd1741: out <= 24'h80d8d7;
        12'd1742: out <= 24'h7ed6e4;
        12'd1743: out <= 24'h7ed6e4;
        12'd1744: out <= 24'h80e20f;
        12'd1745: out <= 24'h82e520;
        12'd1746: out <= 24'h80e32d;
        12'd1747: out <= 24'h7ee13a;
        12'd1748: out <= 24'h81e44c;
        12'd1749: out <= 24'h83e65e;
        12'd1750: out <= 24'h81e46a;
        12'd1751: out <= 24'h80e378;
        12'd1752: out <= 24'h82e689;
        12'd1753: out <= 24'h84e89a;
        12'd1754: out <= 24'h82e6a8;
        12'd1755: out <= 24'h80e5b6;
        12'd1756: out <= 24'h82e8c7;
        12'd1757: out <= 24'h84ead8;
        12'd1758: out <= 24'h82e8e5;
        12'd1759: out <= 24'h82e8e5;
        12'd1760: out <= 24'h80f10c;
        12'd1761: out <= 24'h82f41d;
        12'd1762: out <= 24'h85f62e;
        12'd1763: out <= 24'h83f43c;
        12'd1764: out <= 24'h81f249;
        12'd1765: out <= 24'h83f45a;
        12'd1766: out <= 24'h85f76c;
        12'd1767: out <= 24'h84f679;
        12'd1768: out <= 24'h82f486;
        12'd1769: out <= 24'h84f698;
        12'd1770: out <= 24'h86f9a9;
        12'd1771: out <= 24'h84f8b6;
        12'd1772: out <= 24'h82f6c4;
        12'd1773: out <= 24'h84f8d5;
        12'd1774: out <= 24'h87fbe6;
        12'd1775: out <= 24'h87fbe6;
        12'd1776: out <= 24'h80f10c;
        12'd1777: out <= 24'h82f41d;
        12'd1778: out <= 24'h85f62e;
        12'd1779: out <= 24'h83f43c;
        12'd1780: out <= 24'h81f249;
        12'd1781: out <= 24'h83f45a;
        12'd1782: out <= 24'h85f76c;
        12'd1783: out <= 24'h84f679;
        12'd1784: out <= 24'h82f486;
        12'd1785: out <= 24'h84f698;
        12'd1786: out <= 24'h86f9a9;
        12'd1787: out <= 24'h84f8b6;
        12'd1788: out <= 24'h82f6c4;
        12'd1789: out <= 24'h84f8d5;
        12'd1790: out <= 24'h87fbe6;
        12'd1791: out <= 24'h87fbe6;
        12'd1792: out <= 24'h6a0416;
        12'd1793: out <= 24'h6c0728;
        12'd1794: out <= 24'h6a0635;
        12'd1795: out <= 24'h680442;
        12'd1796: out <= 24'h6b0654;
        12'd1797: out <= 24'h6d0966;
        12'd1798: out <= 24'h6b0872;
        12'd1799: out <= 24'h6a0680;
        12'd1800: out <= 24'h6c0891;
        12'd1801: out <= 24'h6e0ba2;
        12'd1802: out <= 24'h6c09b0;
        12'd1803: out <= 24'h6a07be;
        12'd1804: out <= 24'h6c0acf;
        12'd1805: out <= 24'h6e0ce0;
        12'd1806: out <= 24'h6c0aed;
        12'd1807: out <= 24'h6c0aed;
        12'd1808: out <= 24'h6e1718;
        12'd1809: out <= 24'h6c1624;
        12'd1810: out <= 24'h6a1432;
        12'd1811: out <= 24'h6d1644;
        12'd1812: out <= 24'h701955;
        12'd1813: out <= 24'h6e1862;
        12'd1814: out <= 24'h6c1670;
        12'd1815: out <= 24'h6e1881;
        12'd1816: out <= 24'h701b92;
        12'd1817: out <= 24'h6e1aa0;
        12'd1818: out <= 24'h6c18ad;
        12'd1819: out <= 24'h6e1abe;
        12'd1820: out <= 24'h701cd0;
        12'd1821: out <= 24'h6e1add;
        12'd1822: out <= 24'h6c19ea;
        12'd1823: out <= 24'h6c19ea;
        12'd1824: out <= 24'h732a19;
        12'd1825: out <= 24'h712826;
        12'd1826: out <= 24'h6f2633;
        12'd1827: out <= 24'h722944;
        12'd1828: out <= 24'h742c56;
        12'd1829: out <= 24'h722a64;
        12'd1830: out <= 24'h702871;
        12'd1831: out <= 24'h722b82;
        12'd1832: out <= 24'h742e94;
        12'd1833: out <= 24'h722ca0;
        12'd1834: out <= 24'h702aae;
        12'd1835: out <= 24'h722dc0;
        12'd1836: out <= 24'h7530d1;
        12'd1837: out <= 24'h732ede;
        12'd1838: out <= 24'h712ceb;
        12'd1839: out <= 24'h712ceb;
        12'd1840: out <= 24'h783c1a;
        12'd1841: out <= 24'h763a28;
        12'd1842: out <= 24'h743934;
        12'd1843: out <= 24'h763c46;
        12'd1844: out <= 24'h783e57;
        12'd1845: out <= 24'h763c64;
        12'd1846: out <= 24'h743b72;
        12'd1847: out <= 24'h763e84;
        12'd1848: out <= 24'h784094;
        12'd1849: out <= 24'h763ea2;
        12'd1850: out <= 24'h743daf;
        12'd1851: out <= 24'h723bbc;
        12'd1852: out <= 24'h753ece;
        12'd1853: out <= 24'h7840e0;
        12'd1854: out <= 24'h763eec;
        12'd1855: out <= 24'h763eec;
        12'd1856: out <= 24'h784a17;
        12'd1857: out <= 24'h764924;
        12'd1858: out <= 24'h784c36;
        12'd1859: out <= 24'h7a4e47;
        12'd1860: out <= 24'h784c54;
        12'd1861: out <= 24'h764b62;
        12'd1862: out <= 24'h784e73;
        12'd1863: out <= 24'h7a5084;
        12'd1864: out <= 24'h794e92;
        12'd1865: out <= 24'h774d9e;
        12'd1866: out <= 24'h7950b0;
        12'd1867: out <= 24'h774ebe;
        12'd1868: out <= 24'h754ccb;
        12'd1869: out <= 24'h784edc;
        12'd1870: out <= 24'h7a51ee;
        12'd1871: out <= 24'h7a51ee;
        12'd1872: out <= 24'h785914;
        12'd1873: out <= 24'h7a5c26;
        12'd1874: out <= 24'h7c5e37;
        12'd1875: out <= 24'h7a5c44;
        12'd1876: out <= 24'h785b51;
        12'd1877: out <= 24'h7a5e62;
        12'd1878: out <= 24'h7c6074;
        12'd1879: out <= 24'h7a5e82;
        12'd1880: out <= 24'h795d8e;
        12'd1881: out <= 24'h7c60a0;
        12'd1882: out <= 24'h7e62b2;
        12'd1883: out <= 24'h7c60be;
        12'd1884: out <= 24'h7a5fcc;
        12'd1885: out <= 24'h7c62de;
        12'd1886: out <= 24'h7e64ef;
        12'd1887: out <= 24'h7e64ef;
        12'd1888: out <= 24'h7c6c15;
        12'd1889: out <= 24'h7e6e26;
        12'd1890: out <= 24'h7c6c34;
        12'd1891: out <= 24'h7a6b41;
        12'd1892: out <= 24'h7d6e52;
        12'd1893: out <= 24'h7f7064;
        12'd1894: out <= 24'h7d6e71;
        12'd1895: out <= 24'h7b6d7e;
        12'd1896: out <= 24'h7d7090;
        12'd1897: out <= 24'h8072a2;
        12'd1898: out <= 24'h7e70ae;
        12'd1899: out <= 24'h7c6fbc;
        12'd1900: out <= 24'h7e72cd;
        12'd1901: out <= 24'h8074de;
        12'd1902: out <= 24'h7e72ec;
        12'd1903: out <= 24'h7e72ec;
        12'd1904: out <= 24'h807e16;
        12'd1905: out <= 24'h7e7c24;
        12'd1906: out <= 24'h7c7b31;
        12'd1907: out <= 24'h7e7e42;
        12'd1908: out <= 24'h818054;
        12'd1909: out <= 24'h807e60;
        12'd1910: out <= 24'h7e7d6e;
        12'd1911: out <= 24'h808080;
        12'd1912: out <= 24'h828291;
        12'd1913: out <= 24'h80809e;
        12'd1914: out <= 24'h7e7fac;
        12'd1915: out <= 24'h8082bc;
        12'd1916: out <= 24'h8284ce;
        12'd1917: out <= 24'h8082dc;
        12'd1918: out <= 24'h7e80e9;
        12'd1919: out <= 24'h7e80e9;
        12'd1920: out <= 24'h818d13;
        12'd1921: out <= 24'h7f8b20;
        12'd1922: out <= 24'h818e32;
        12'd1923: out <= 24'h839044;
        12'd1924: out <= 24'h818e50;
        12'd1925: out <= 24'h808d5e;
        12'd1926: out <= 24'h82906f;
        12'd1927: out <= 24'h849280;
        12'd1928: out <= 24'h82908e;
        12'd1929: out <= 24'h808f9c;
        12'd1930: out <= 24'h8292ad;
        12'd1931: out <= 24'h8494be;
        12'd1932: out <= 24'h8392cb;
        12'd1933: out <= 24'h8191d8;
        12'd1934: out <= 24'h8394ea;
        12'd1935: out <= 24'h8394ea;
        12'd1936: out <= 24'h819b10;
        12'd1937: out <= 24'h849e22;
        12'd1938: out <= 24'h86a033;
        12'd1939: out <= 24'h849e40;
        12'd1940: out <= 24'h829d4e;
        12'd1941: out <= 24'h84a05f;
        12'd1942: out <= 24'h86a270;
        12'd1943: out <= 24'h84a07e;
        12'd1944: out <= 24'h829f8b;
        12'd1945: out <= 24'h84a29c;
        12'd1946: out <= 24'h86a4ae;
        12'd1947: out <= 24'h84a2bb;
        12'd1948: out <= 24'h83a1c8;
        12'd1949: out <= 24'h86a4da;
        12'd1950: out <= 24'h88a6eb;
        12'd1951: out <= 24'h88a6eb;
        12'd1952: out <= 24'h85ae11;
        12'd1953: out <= 24'h88b022;
        12'd1954: out <= 24'h8ab334;
        12'd1955: out <= 24'h88b242;
        12'd1956: out <= 24'h86b04f;
        12'd1957: out <= 24'h88b260;
        12'd1958: out <= 24'h8ab472;
        12'd1959: out <= 24'h88b37e;
        12'd1960: out <= 24'h87b28c;
        12'd1961: out <= 24'h89b49e;
        12'd1962: out <= 24'h87b2ab;
        12'd1963: out <= 24'h85b1b8;
        12'd1964: out <= 24'h87b4c9;
        12'd1965: out <= 24'h8ab6da;
        12'd1966: out <= 24'h88b4e8;
        12'd1967: out <= 24'h88b4e8;
        12'd1968: out <= 24'h8ac112;
        12'd1969: out <= 24'h88bf20;
        12'd1970: out <= 24'h8ac231;
        12'd1971: out <= 24'h8cc442;
        12'd1972: out <= 24'h8ac250;
        12'd1973: out <= 24'h88c05e;
        12'd1974: out <= 24'h8ac36e;
        12'd1975: out <= 24'h8cc680;
        12'd1976: out <= 24'h8bc48d;
        12'd1977: out <= 24'h89c29a;
        12'd1978: out <= 24'h87c1a8;
        12'd1979: out <= 24'h8ac4ba;
        12'd1980: out <= 24'h8cc6ca;
        12'd1981: out <= 24'h8ac4d8;
        12'd1982: out <= 24'h88c3e5;
        12'd1983: out <= 24'h88c3e5;
        12'd1984: out <= 24'h8ed414;
        12'd1985: out <= 24'h8cd221;
        12'd1986: out <= 24'h8ad02e;
        12'd1987: out <= 24'h8cd240;
        12'd1988: out <= 24'h8fd451;
        12'd1989: out <= 24'h8dd35e;
        12'd1990: out <= 24'h8bd26c;
        12'd1991: out <= 24'h8dd47c;
        12'd1992: out <= 24'h8fd68e;
        12'd1993: out <= 24'h8dd59c;
        12'd1994: out <= 24'h8bd4a9;
        12'd1995: out <= 24'h8ed6ba;
        12'd1996: out <= 24'h90d8cc;
        12'd1997: out <= 24'h8ed7d9;
        12'd1998: out <= 24'h8cd6e6;
        12'd1999: out <= 24'h8cd6e6;
        12'd2000: out <= 24'h92e615;
        12'd2001: out <= 24'h90e422;
        12'd2002: out <= 24'h8ee22f;
        12'd2003: out <= 24'h90e540;
        12'd2004: out <= 24'h93e852;
        12'd2005: out <= 24'h91e660;
        12'd2006: out <= 24'h8fe46c;
        12'd2007: out <= 24'h92e67e;
        12'd2008: out <= 24'h94e990;
        12'd2009: out <= 24'h92e89c;
        12'd2010: out <= 24'h90e6aa;
        12'd2011: out <= 24'h92e8bc;
        12'd2012: out <= 24'h94ebcd;
        12'd2013: out <= 24'h92eada;
        12'd2014: out <= 24'h90e8e8;
        12'd2015: out <= 24'h90e8e8;
        12'd2016: out <= 24'h92f412;
        12'd2017: out <= 24'h90f31f;
        12'd2018: out <= 24'h93f630;
        12'd2019: out <= 24'h95f842;
        12'd2020: out <= 24'h93f64f;
        12'd2021: out <= 24'h91f45c;
        12'd2022: out <= 24'h93f66e;
        12'd2023: out <= 24'h96f980;
        12'd2024: out <= 24'h94f88c;
        12'd2025: out <= 24'h92f69a;
        12'd2026: out <= 24'h94f8ab;
        12'd2027: out <= 24'h96fbbc;
        12'd2028: out <= 24'h94faca;
        12'd2029: out <= 24'h92f8d8;
        12'd2030: out <= 24'h95fae8;
        12'd2031: out <= 24'h95fae8;
        12'd2032: out <= 24'h92f412;
        12'd2033: out <= 24'h90f31f;
        12'd2034: out <= 24'h93f630;
        12'd2035: out <= 24'h95f842;
        12'd2036: out <= 24'h93f64f;
        12'd2037: out <= 24'h91f45c;
        12'd2038: out <= 24'h93f66e;
        12'd2039: out <= 24'h96f980;
        12'd2040: out <= 24'h94f88c;
        12'd2041: out <= 24'h92f69a;
        12'd2042: out <= 24'h94f8ab;
        12'd2043: out <= 24'h96fbbc;
        12'd2044: out <= 24'h94faca;
        12'd2045: out <= 24'h92f8d8;
        12'd2046: out <= 24'h95fae8;
        12'd2047: out <= 24'h95fae8;
        12'd2048: out <= 24'h780419;
        12'd2049: out <= 24'h7a062a;
        12'd2050: out <= 24'h7d093b;
        12'd2051: out <= 24'h7b0848;
        12'd2052: out <= 24'h790656;
        12'd2053: out <= 24'h7b0868;
        12'd2054: out <= 24'h7d0b79;
        12'd2055: out <= 24'h7c0a86;
        12'd2056: out <= 24'h7a0893;
        12'd2057: out <= 24'h7c0aa4;
        12'd2058: out <= 24'h7e0db6;
        12'd2059: out <= 24'h7c0bc4;
        12'd2060: out <= 24'h7a09d1;
        12'd2061: out <= 24'h7c0ce2;
        12'd2062: out <= 24'h7f0ef3;
        12'd2063: out <= 24'h7f0ef3;
        12'd2064: out <= 24'h7c161a;
        12'd2065: out <= 24'h7a1527;
        12'd2066: out <= 24'h7d1838;
        12'd2067: out <= 24'h801a4a;
        12'd2068: out <= 24'h7e1857;
        12'd2069: out <= 24'h7c1764;
        12'd2070: out <= 24'h7e1a76;
        12'd2071: out <= 24'h801c88;
        12'd2072: out <= 24'h7e1a94;
        12'd2073: out <= 24'h7c19a2;
        12'd2074: out <= 24'h7e1cb3;
        12'd2075: out <= 24'h801ec4;
        12'd2076: out <= 24'h7e1cd2;
        12'd2077: out <= 24'h7c1adf;
        12'd2078: out <= 24'h7f1cf0;
        12'd2079: out <= 24'h7f1cf0;
        12'd2080: out <= 24'h81291b;
        12'd2081: out <= 24'h7f2828;
        12'd2082: out <= 24'h7d2635;
        12'd2083: out <= 24'h802846;
        12'd2084: out <= 24'h822b58;
        12'd2085: out <= 24'h802a66;
        12'd2086: out <= 24'h7e2873;
        12'd2087: out <= 24'h802a84;
        12'd2088: out <= 24'h822d96;
        12'd2089: out <= 24'h802ca3;
        12'd2090: out <= 24'h7e2ab0;
        12'd2091: out <= 24'h802cc2;
        12'd2092: out <= 24'h832fd3;
        12'd2093: out <= 24'h812de0;
        12'd2094: out <= 24'h7f2bed;
        12'd2095: out <= 24'h7f2bed;
        12'd2096: out <= 24'h863c1c;
        12'd2097: out <= 24'h843a2a;
        12'd2098: out <= 24'h823836;
        12'd2099: out <= 24'h843b48;
        12'd2100: out <= 24'h863e59;
        12'd2101: out <= 24'h843c66;
        12'd2102: out <= 24'h823a74;
        12'd2103: out <= 24'h843d86;
        12'd2104: out <= 24'h864097;
        12'd2105: out <= 24'h843ea4;
        12'd2106: out <= 24'h823cb1;
        12'd2107: out <= 24'h803abe;
        12'd2108: out <= 24'h833dd0;
        12'd2109: out <= 24'h8640e2;
        12'd2110: out <= 24'h843eee;
        12'd2111: out <= 24'h843eee;
        12'd2112: out <= 24'h8a4e1d;
        12'd2113: out <= 24'h884c2a;
        12'd2114: out <= 24'h864b38;
        12'd2115: out <= 24'h884e49;
        12'd2116: out <= 24'h8a505a;
        12'd2117: out <= 24'h884e68;
        12'd2118: out <= 24'h864d75;
        12'd2119: out <= 24'h885086;
        12'd2120: out <= 24'h8b5298;
        12'd2121: out <= 24'h8950a5;
        12'd2122: out <= 24'h874fb2;
        12'd2123: out <= 24'h854dc0;
        12'd2124: out <= 24'h834bcd;
        12'd2125: out <= 24'h864ede;
        12'd2126: out <= 24'h8850f0;
        12'd2127: out <= 24'h8850f0;
        12'd2128: out <= 24'h8a5c1a;
        12'd2129: out <= 24'h8c5f2c;
        12'd2130: out <= 24'h8a5e39;
        12'd2131: out <= 24'h885c46;
        12'd2132: out <= 24'h8a5e57;
        12'd2133: out <= 24'h8c6168;
        12'd2134: out <= 24'h8a6076;
        12'd2135: out <= 24'h885e84;
        12'd2136: out <= 24'h8b6095;
        12'd2137: out <= 24'h8e63a6;
        12'd2138: out <= 24'h8c62b4;
        12'd2139: out <= 24'h8a60c0;
        12'd2140: out <= 24'h885ece;
        12'd2141: out <= 24'h8a60e0;
        12'd2142: out <= 24'h8c63f1;
        12'd2143: out <= 24'h8c63f1;
        12'd2144: out <= 24'h8a6b17;
        12'd2145: out <= 24'h8c6e28;
        12'd2146: out <= 24'h8e703a;
        12'd2147: out <= 24'h8c6e47;
        12'd2148: out <= 24'h8b6d54;
        12'd2149: out <= 24'h8d7066;
        12'd2150: out <= 24'h8f7277;
        12'd2151: out <= 24'h8d7084;
        12'd2152: out <= 24'h8b6f92;
        12'd2153: out <= 24'h8e72a4;
        12'd2154: out <= 24'h9074b5;
        12'd2155: out <= 24'h8e72c2;
        12'd2156: out <= 24'h8c71cf;
        12'd2157: out <= 24'h8e74e0;
        12'd2158: out <= 24'h9076f2;
        12'd2159: out <= 24'h9076f2;
        12'd2160: out <= 24'h8e7e18;
        12'd2161: out <= 24'h8c7c26;
        12'd2162: out <= 24'h8e7e37;
        12'd2163: out <= 24'h908148;
        12'd2164: out <= 24'h8f8056;
        12'd2165: out <= 24'h8e7e62;
        12'd2166: out <= 24'h908074;
        12'd2167: out <= 24'h928386;
        12'd2168: out <= 24'h908293;
        12'd2169: out <= 24'h8e80a0;
        12'd2170: out <= 24'h9082b2;
        12'd2171: out <= 24'h9285c3;
        12'd2172: out <= 24'h9084d0;
        12'd2173: out <= 24'h8e82de;
        12'd2174: out <= 24'h9084ef;
        12'd2175: out <= 24'h9084ef;
        12'd2176: out <= 24'h939119;
        12'd2177: out <= 24'h918f26;
        12'd2178: out <= 24'h8f8d34;
        12'd2179: out <= 24'h919046;
        12'd2180: out <= 24'h939257;
        12'd2181: out <= 24'h929064;
        12'd2182: out <= 24'h908f71;
        12'd2183: out <= 24'h929282;
        12'd2184: out <= 24'h949494;
        12'd2185: out <= 24'h9292a2;
        12'd2186: out <= 24'h9091af;
        12'd2187: out <= 24'h9294c0;
        12'd2188: out <= 24'h9596d1;
        12'd2189: out <= 24'h9394de;
        12'd2190: out <= 24'h9193ec;
        12'd2191: out <= 24'h9193ec;
        12'd2192: out <= 24'h939f16;
        12'd2193: out <= 24'h96a228;
        12'd2194: out <= 24'h94a035;
        12'd2195: out <= 24'h929e42;
        12'd2196: out <= 24'h94a054;
        12'd2197: out <= 24'h96a366;
        12'd2198: out <= 24'h94a272;
        12'd2199: out <= 24'h92a080;
        12'd2200: out <= 24'h94a291;
        12'd2201: out <= 24'h96a5a2;
        12'd2202: out <= 24'h94a4b0;
        12'd2203: out <= 24'h92a2bd;
        12'd2204: out <= 24'h95a4ce;
        12'd2205: out <= 24'h98a7e0;
        12'd2206: out <= 24'h96a6ed;
        12'd2207: out <= 24'h96a6ed;
        12'd2208: out <= 24'h93ad13;
        12'd2209: out <= 24'h96b024;
        12'd2210: out <= 24'h98b236;
        12'd2211: out <= 24'h96b044;
        12'd2212: out <= 24'h94af51;
        12'd2213: out <= 24'h96b262;
        12'd2214: out <= 24'h98b474;
        12'd2215: out <= 24'h96b281;
        12'd2216: out <= 24'h95b18e;
        12'd2217: out <= 24'h97b4a0;
        12'd2218: out <= 24'h99b6b1;
        12'd2219: out <= 24'h97b4be;
        12'd2220: out <= 24'h95b3cb;
        12'd2221: out <= 24'h98b6dc;
        12'd2222: out <= 24'h9ab8ee;
        12'd2223: out <= 24'h9ab8ee;
        12'd2224: out <= 24'h98c014;
        12'd2225: out <= 24'h96be22;
        12'd2226: out <= 24'h98c033;
        12'd2227: out <= 24'h9ac344;
        12'd2228: out <= 24'h98c252;
        12'd2229: out <= 24'h96c060;
        12'd2230: out <= 24'h98c271;
        12'd2231: out <= 24'h9ac582;
        12'd2232: out <= 24'h99c48f;
        12'd2233: out <= 24'h97c29c;
        12'd2234: out <= 24'h99c4ae;
        12'd2235: out <= 24'h9cc7c0;
        12'd2236: out <= 24'h9ac6cc;
        12'd2237: out <= 24'h98c4da;
        12'd2238: out <= 24'h9ac6eb;
        12'd2239: out <= 24'h9ac6eb;
        12'd2240: out <= 24'h9cd316;
        12'd2241: out <= 24'h9ad123;
        12'd2242: out <= 24'h98cf30;
        12'd2243: out <= 24'h9ad242;
        12'd2244: out <= 24'h9dd453;
        12'd2245: out <= 24'h9bd260;
        12'd2246: out <= 24'h99d16e;
        12'd2247: out <= 24'h9bd47f;
        12'd2248: out <= 24'h9dd690;
        12'd2249: out <= 24'h9bd49e;
        12'd2250: out <= 24'h99d3ab;
        12'd2251: out <= 24'h9cd6bc;
        12'd2252: out <= 24'h9ed8ce;
        12'd2253: out <= 24'h9cd6db;
        12'd2254: out <= 24'h9ad5e8;
        12'd2255: out <= 24'h9ad5e8;
        12'd2256: out <= 24'ha0e617;
        12'd2257: out <= 24'h9ee424;
        12'd2258: out <= 24'h9ce231;
        12'd2259: out <= 24'h9ee442;
        12'd2260: out <= 24'ha1e754;
        12'd2261: out <= 24'h9fe562;
        12'd2262: out <= 24'h9de46f;
        12'd2263: out <= 24'ha0e680;
        12'd2264: out <= 24'ha2e892;
        12'd2265: out <= 24'ha0e79e;
        12'd2266: out <= 24'h9ee6ac;
        12'd2267: out <= 24'ha0e8be;
        12'd2268: out <= 24'ha2eacf;
        12'd2269: out <= 24'ha0e9dc;
        12'd2270: out <= 24'h9ee8ea;
        12'd2271: out <= 24'h9ee8ea;
        12'd2272: out <= 24'ha5f818;
        12'd2273: out <= 24'ha3f625;
        12'd2274: out <= 24'ha1f532;
        12'd2275: out <= 24'ha3f844;
        12'd2276: out <= 24'ha5fa55;
        12'd2277: out <= 24'ha3f862;
        12'd2278: out <= 24'ha1f670;
        12'd2279: out <= 24'ha4f882;
        12'd2280: out <= 24'ha6fb93;
        12'd2281: out <= 24'ha4faa0;
        12'd2282: out <= 24'ha2f8ad;
        12'd2283: out <= 24'ha4fabe;
        12'd2284: out <= 24'ha7fdd0;
        12'd2285: out <= 24'ha5fcde;
        12'd2286: out <= 24'ha3faeb;
        12'd2287: out <= 24'ha3faeb;
        12'd2288: out <= 24'ha5f818;
        12'd2289: out <= 24'ha3f625;
        12'd2290: out <= 24'ha1f532;
        12'd2291: out <= 24'ha3f844;
        12'd2292: out <= 24'ha5fa55;
        12'd2293: out <= 24'ha3f862;
        12'd2294: out <= 24'ha1f670;
        12'd2295: out <= 24'ha4f882;
        12'd2296: out <= 24'ha6fb93;
        12'd2297: out <= 24'ha4faa0;
        12'd2298: out <= 24'ha2f8ad;
        12'd2299: out <= 24'ha4fabe;
        12'd2300: out <= 24'ha7fdd0;
        12'd2301: out <= 24'ha5fcde;
        12'd2302: out <= 24'ha3faeb;
        12'd2303: out <= 24'ha3faeb;
        12'd2304: out <= 24'h8a081f;
        12'd2305: out <= 24'h88062c;
        12'd2306: out <= 24'h8b083d;
        12'd2307: out <= 24'h8d0b4e;
        12'd2308: out <= 24'h8b0a5c;
        12'd2309: out <= 24'h89086a;
        12'd2310: out <= 24'h8b0a7b;
        12'd2311: out <= 24'h8e0d8c;
        12'd2312: out <= 24'h8c0c9a;
        12'd2313: out <= 24'h8a0aa6;
        12'd2314: out <= 24'h8c0cb8;
        12'd2315: out <= 24'h8e0fca;
        12'd2316: out <= 24'h8c0dd7;
        12'd2317: out <= 24'h8a0be4;
        12'd2318: out <= 24'h8d0ef5;
        12'd2319: out <= 24'h8d0ef5;
        12'd2320: out <= 24'h8a161c;
        12'd2321: out <= 24'h8c182e;
        12'd2322: out <= 24'h8f1b3e;
        12'd2323: out <= 24'h8e1a4c;
        12'd2324: out <= 24'h8c1859;
        12'd2325: out <= 24'h8e1a6a;
        12'd2326: out <= 24'h901d7c;
        12'd2327: out <= 24'h8e1c8a;
        12'd2328: out <= 24'h8c1a96;
        12'd2329: out <= 24'h8e1ca8;
        12'd2330: out <= 24'h901fb9;
        12'd2331: out <= 24'h8e1dc6;
        12'd2332: out <= 24'h8c1bd4;
        12'd2333: out <= 24'h8e1ee6;
        12'd2334: out <= 24'h9120f6;
        12'd2335: out <= 24'h9120f6;
        12'd2336: out <= 24'h8f281d;
        12'd2337: out <= 24'h912b2e;
        12'd2338: out <= 24'h8f2a3c;
        12'd2339: out <= 24'h8e2848;
        12'd2340: out <= 24'h902a5a;
        12'd2341: out <= 24'h922d6c;
        12'd2342: out <= 24'h902c79;
        12'd2343: out <= 24'h8e2a86;
        12'd2344: out <= 24'h902c98;
        12'd2345: out <= 24'h922fa9;
        12'd2346: out <= 24'h902eb6;
        12'd2347: out <= 24'h8e2cc4;
        12'd2348: out <= 24'h912ed5;
        12'd2349: out <= 24'h9330e6;
        12'd2350: out <= 24'h912ef4;
        12'd2351: out <= 24'h912ef4;
        12'd2352: out <= 24'h943b1e;
        12'd2353: out <= 24'h923a2c;
        12'd2354: out <= 24'h903838;
        12'd2355: out <= 24'h923a4a;
        12'd2356: out <= 24'h943d5c;
        12'd2357: out <= 24'h923c68;
        12'd2358: out <= 24'h903a76;
        12'd2359: out <= 24'h923c88;
        12'd2360: out <= 24'h943f99;
        12'd2361: out <= 24'h923ea6;
        12'd2362: out <= 24'h903cb3;
        12'd2363: out <= 24'h933ec4;
        12'd2364: out <= 24'h9641d6;
        12'd2365: out <= 24'h943fe4;
        12'd2366: out <= 24'h923df0;
        12'd2367: out <= 24'h923df0;
        12'd2368: out <= 24'h984e1f;
        12'd2369: out <= 24'h964c2c;
        12'd2370: out <= 24'h944a3a;
        12'd2371: out <= 24'h964d4c;
        12'd2372: out <= 24'h98505c;
        12'd2373: out <= 24'h964e6a;
        12'd2374: out <= 24'h944c77;
        12'd2375: out <= 24'h964f88;
        12'd2376: out <= 24'h99529a;
        12'd2377: out <= 24'h9750a7;
        12'd2378: out <= 24'h954eb4;
        12'd2379: out <= 24'h9851c6;
        12'd2380: out <= 24'h964fd3;
        12'd2381: out <= 24'h944de0;
        12'd2382: out <= 24'h9650f2;
        12'd2383: out <= 24'h9650f2;
        12'd2384: out <= 24'h985c1c;
        12'd2385: out <= 24'h9a5e2e;
        12'd2386: out <= 24'h985d3b;
        12'd2387: out <= 24'h965c48;
        12'd2388: out <= 24'h985e5a;
        12'd2389: out <= 24'h9a606a;
        12'd2390: out <= 24'h985f78;
        12'd2391: out <= 24'h965e86;
        12'd2392: out <= 24'h996097;
        12'd2393: out <= 24'h9c62a8;
        12'd2394: out <= 24'h9a61b6;
        12'd2395: out <= 24'h9860c2;
        12'd2396: out <= 24'h965ed0;
        12'd2397: out <= 24'h9860e2;
        12'd2398: out <= 24'h9a62f3;
        12'd2399: out <= 24'h9a62f3;
        12'd2400: out <= 24'h986a19;
        12'd2401: out <= 24'h9a6d2a;
        12'd2402: out <= 24'h9c703c;
        12'd2403: out <= 24'h9a6e4a;
        12'd2404: out <= 24'h996c56;
        12'd2405: out <= 24'h9b6f68;
        12'd2406: out <= 24'h9d7279;
        12'd2407: out <= 24'h9b7086;
        12'd2408: out <= 24'h996e94;
        12'd2409: out <= 24'h9c71a6;
        12'd2410: out <= 24'h9e74b7;
        12'd2411: out <= 24'h9c72c4;
        12'd2412: out <= 24'h9a70d1;
        12'd2413: out <= 24'h9c73e2;
        12'd2414: out <= 24'h9e76f4;
        12'd2415: out <= 24'h9e76f4;
        12'd2416: out <= 24'h9c7d1a;
        12'd2417: out <= 24'h9e802c;
        12'd2418: out <= 24'ha0823d;
        12'd2419: out <= 24'h9e804a;
        12'd2420: out <= 24'h9d7f58;
        12'd2421: out <= 24'ha08269;
        12'd2422: out <= 24'ha2847a;
        12'd2423: out <= 24'ha08288;
        12'd2424: out <= 24'h9e8195;
        12'd2425: out <= 24'ha084a6;
        12'd2426: out <= 24'ha286b8;
        12'd2427: out <= 24'ha084c5;
        12'd2428: out <= 24'h9e83d2;
        12'd2429: out <= 24'ha086e4;
        12'd2430: out <= 24'ha288f5;
        12'd2431: out <= 24'ha288f5;
        12'd2432: out <= 24'ha1901b;
        12'd2433: out <= 24'ha3922c;
        12'd2434: out <= 24'ha1903a;
        12'd2435: out <= 24'h9f8f48;
        12'd2436: out <= 24'ha19259;
        12'd2437: out <= 24'ha4946a;
        12'd2438: out <= 24'ha29278;
        12'd2439: out <= 24'ha09184;
        12'd2440: out <= 24'ha29496;
        12'd2441: out <= 24'ha496a8;
        12'd2442: out <= 24'ha294b5;
        12'd2443: out <= 24'ha093c2;
        12'd2444: out <= 24'ha396d3;
        12'd2445: out <= 24'ha598e4;
        12'd2446: out <= 24'ha396f2;
        12'd2447: out <= 24'ha396f2;
        12'd2448: out <= 24'ha5a31c;
        12'd2449: out <= 24'ha4a12a;
        12'd2450: out <= 24'ha29f37;
        12'd2451: out <= 24'ha4a248;
        12'd2452: out <= 24'ha6a45a;
        12'd2453: out <= 24'ha4a268;
        12'd2454: out <= 24'ha2a174;
        12'd2455: out <= 24'ha4a486;
        12'd2456: out <= 24'ha6a697;
        12'd2457: out <= 24'ha4a4a4;
        12'd2458: out <= 24'ha2a3b2;
        12'd2459: out <= 24'ha4a6c4;
        12'd2460: out <= 24'ha7a8d4;
        12'd2461: out <= 24'ha6a6e2;
        12'd2462: out <= 24'ha4a5ef;
        12'd2463: out <= 24'ha4a5ef;
        12'd2464: out <= 24'ha5b11a;
        12'd2465: out <= 24'ha4af26;
        12'd2466: out <= 24'ha6b238;
        12'd2467: out <= 24'ha8b44a;
        12'd2468: out <= 24'ha6b257;
        12'd2469: out <= 24'ha4b164;
        12'd2470: out <= 24'ha6b476;
        12'd2471: out <= 24'ha8b687;
        12'd2472: out <= 24'ha7b494;
        12'd2473: out <= 24'ha5b3a2;
        12'd2474: out <= 24'ha7b6b3;
        12'd2475: out <= 24'ha9b8c4;
        12'd2476: out <= 24'ha7b6d2;
        12'd2477: out <= 24'ha6b5de;
        12'd2478: out <= 24'ha8b8f0;
        12'd2479: out <= 24'ha8b8f0;
        12'd2480: out <= 24'ha6c016;
        12'd2481: out <= 24'ha8c228;
        12'd2482: out <= 24'haac43a;
        12'd2483: out <= 24'ha8c246;
        12'd2484: out <= 24'ha6c154;
        12'd2485: out <= 24'ha8c466;
        12'd2486: out <= 24'haac677;
        12'd2487: out <= 24'ha8c484;
        12'd2488: out <= 24'ha7c391;
        12'd2489: out <= 24'haac6a2;
        12'd2490: out <= 24'hacc8b4;
        12'd2491: out <= 24'haac6c2;
        12'd2492: out <= 24'ha8c5ce;
        12'd2493: out <= 24'haac8e0;
        12'd2494: out <= 24'haccaf2;
        12'd2495: out <= 24'haccaf2;
        12'd2496: out <= 24'haad218;
        12'd2497: out <= 24'hacd52a;
        12'd2498: out <= 24'haad336;
        12'd2499: out <= 24'ha8d144;
        12'd2500: out <= 24'habd455;
        12'd2501: out <= 24'hadd666;
        12'd2502: out <= 24'habd474;
        12'd2503: out <= 24'ha9d381;
        12'd2504: out <= 24'habd692;
        12'd2505: out <= 24'haed8a4;
        12'd2506: out <= 24'hacd6b1;
        12'd2507: out <= 24'haad5be;
        12'd2508: out <= 24'hacd8d0;
        12'd2509: out <= 24'haedae2;
        12'd2510: out <= 24'hacd8ee;
        12'd2511: out <= 24'hacd8ee;
        12'd2512: out <= 24'haee519;
        12'd2513: out <= 24'hace426;
        12'd2514: out <= 24'haae234;
        12'd2515: out <= 24'hace444;
        12'd2516: out <= 24'hafe656;
        12'd2517: out <= 24'hade464;
        12'd2518: out <= 24'habe371;
        12'd2519: out <= 24'haee682;
        12'd2520: out <= 24'hb0e894;
        12'd2521: out <= 24'haee6a0;
        12'd2522: out <= 24'hace5ae;
        12'd2523: out <= 24'haee8c0;
        12'd2524: out <= 24'hb0ead1;
        12'd2525: out <= 24'haee8de;
        12'd2526: out <= 24'hace7ec;
        12'd2527: out <= 24'hace7ec;
        12'd2528: out <= 24'hb3f81a;
        12'd2529: out <= 24'hb1f628;
        12'd2530: out <= 24'haff434;
        12'd2531: out <= 24'hb1f746;
        12'd2532: out <= 24'hb3fa57;
        12'd2533: out <= 24'hb1f864;
        12'd2534: out <= 24'haff672;
        12'd2535: out <= 24'hb2f884;
        12'd2536: out <= 24'hb4fa95;
        12'd2537: out <= 24'hb2f9a2;
        12'd2538: out <= 24'hb0f8af;
        12'd2539: out <= 24'hb2fac0;
        12'd2540: out <= 24'hb5fcd2;
        12'd2541: out <= 24'hb3fbe0;
        12'd2542: out <= 24'hb1faed;
        12'd2543: out <= 24'hb1faed;
        12'd2544: out <= 24'hb3f81a;
        12'd2545: out <= 24'hb1f628;
        12'd2546: out <= 24'haff434;
        12'd2547: out <= 24'hb1f746;
        12'd2548: out <= 24'hb3fa57;
        12'd2549: out <= 24'hb1f864;
        12'd2550: out <= 24'haff672;
        12'd2551: out <= 24'hb2f884;
        12'd2552: out <= 24'hb4fa95;
        12'd2553: out <= 24'hb2f9a2;
        12'd2554: out <= 24'hb0f8af;
        12'd2555: out <= 24'hb2fac0;
        12'd2556: out <= 24'hb5fcd2;
        12'd2557: out <= 24'hb3fbe0;
        12'd2558: out <= 24'hb1faed;
        12'd2559: out <= 24'hb1faed;
        12'd2560: out <= 24'h9c0b25;
        12'd2561: out <= 24'h9a0a32;
        12'd2562: out <= 24'h99083f;
        12'd2563: out <= 24'h9b0a50;
        12'd2564: out <= 24'h9d0d62;
        12'd2565: out <= 24'h9b0c70;
        12'd2566: out <= 24'h990a7d;
        12'd2567: out <= 24'h9c0c8e;
        12'd2568: out <= 24'h9e0fa0;
        12'd2569: out <= 24'h9c0ead;
        12'd2570: out <= 24'h9a0cba;
        12'd2571: out <= 24'h9c0ecc;
        12'd2572: out <= 24'h9e11dd;
        12'd2573: out <= 24'h9c0fea;
        12'd2574: out <= 24'h9b0df7;
        12'd2575: out <= 24'h9b0df7;
        12'd2576: out <= 24'h9c1a22;
        12'd2577: out <= 24'h9e1c34;
        12'd2578: out <= 24'h9d1a40;
        12'd2579: out <= 24'h9c194e;
        12'd2580: out <= 24'h9e1c5f;
        12'd2581: out <= 24'ha01e70;
        12'd2582: out <= 24'h9e1c7e;
        12'd2583: out <= 24'h9c1b8c;
        12'd2584: out <= 24'h9e1e9d;
        12'd2585: out <= 24'ha020ae;
        12'd2586: out <= 24'h9e1ebb;
        12'd2587: out <= 24'h9c1cc8;
        12'd2588: out <= 24'h9e1fda;
        12'd2589: out <= 24'ha022ec;
        12'd2590: out <= 24'h9f20f8;
        12'd2591: out <= 24'h9f20f8;
        12'd2592: out <= 24'h9d281f;
        12'd2593: out <= 24'h9f2a30;
        12'd2594: out <= 24'ha12d42;
        12'd2595: out <= 24'ha02c4f;
        12'd2596: out <= 24'h9e2a5c;
        12'd2597: out <= 24'ha02c6e;
        12'd2598: out <= 24'ha22f7f;
        12'd2599: out <= 24'ha02e8c;
        12'd2600: out <= 24'h9e2c9a;
        12'd2601: out <= 24'ha02eab;
        12'd2602: out <= 24'ha331bc;
        12'd2603: out <= 24'ha12fca;
        12'd2604: out <= 24'h9f2dd7;
        12'd2605: out <= 24'ha130e8;
        12'd2606: out <= 24'ha332fa;
        12'd2607: out <= 24'ha332fa;
        12'd2608: out <= 24'ha23a20;
        12'd2609: out <= 24'ha0392e;
        12'd2610: out <= 24'ha23c3f;
        12'd2611: out <= 24'ha43e50;
        12'd2612: out <= 24'ha23c5e;
        12'd2613: out <= 24'ha03b6a;
        12'd2614: out <= 24'ha23e7c;
        12'd2615: out <= 24'ha4408e;
        12'd2616: out <= 24'ha23e9b;
        12'd2617: out <= 24'ha03da8;
        12'd2618: out <= 24'ha340b9;
        12'd2619: out <= 24'ha642ca;
        12'd2620: out <= 24'ha440d8;
        12'd2621: out <= 24'ha23ee6;
        12'd2622: out <= 24'ha440f7;
        12'd2623: out <= 24'ha440f7;
        12'd2624: out <= 24'ha64d21;
        12'd2625: out <= 24'ha44c2e;
        12'd2626: out <= 24'ha24a3c;
        12'd2627: out <= 24'ha44c4e;
        12'd2628: out <= 24'ha64f5f;
        12'd2629: out <= 24'ha44e6c;
        12'd2630: out <= 24'ha24c79;
        12'd2631: out <= 24'ha44e8a;
        12'd2632: out <= 24'ha7519c;
        12'd2633: out <= 24'ha550a9;
        12'd2634: out <= 24'ha34eb6;
        12'd2635: out <= 24'ha650c8;
        12'd2636: out <= 24'ha853d9;
        12'd2637: out <= 24'ha651e6;
        12'd2638: out <= 24'ha44ff4;
        12'd2639: out <= 24'ha44ff4;
        12'd2640: out <= 24'ha65c1e;
        12'd2641: out <= 24'ha85e30;
        12'd2642: out <= 24'ha65c3d;
        12'd2643: out <= 24'ha45b4a;
        12'd2644: out <= 24'ha65e5c;
        12'd2645: out <= 24'ha8606d;
        12'd2646: out <= 24'ha65e7a;
        12'd2647: out <= 24'ha45d88;
        12'd2648: out <= 24'ha76099;
        12'd2649: out <= 24'haa62aa;
        12'd2650: out <= 24'ha860b8;
        12'd2651: out <= 24'ha65fc4;
        12'd2652: out <= 24'ha862d6;
        12'd2653: out <= 24'haa64e8;
        12'd2654: out <= 24'ha862f5;
        12'd2655: out <= 24'ha862f5;
        12'd2656: out <= 24'ha66a1b;
        12'd2657: out <= 24'ha86c2c;
        12'd2658: out <= 24'haa6f3e;
        12'd2659: out <= 24'ha86e4c;
        12'd2660: out <= 24'ha76c59;
        12'd2661: out <= 24'ha96e6a;
        12'd2662: out <= 24'hab717b;
        12'd2663: out <= 24'ha97088;
        12'd2664: out <= 24'ha76e96;
        12'd2665: out <= 24'haa70a8;
        12'd2666: out <= 24'hac73b9;
        12'd2667: out <= 24'haa72c6;
        12'd2668: out <= 24'ha870d3;
        12'd2669: out <= 24'haa72e4;
        12'd2670: out <= 24'hac75f6;
        12'd2671: out <= 24'hac75f6;
        12'd2672: out <= 24'haa7c1c;
        12'd2673: out <= 24'hac7f2e;
        12'd2674: out <= 24'hae823f;
        12'd2675: out <= 24'hac804c;
        12'd2676: out <= 24'hab7e5a;
        12'd2677: out <= 24'hae816c;
        12'd2678: out <= 24'hb0847c;
        12'd2679: out <= 24'hae828a;
        12'd2680: out <= 24'hac8097;
        12'd2681: out <= 24'hae83a8;
        12'd2682: out <= 24'hb086ba;
        12'd2683: out <= 24'hae84c7;
        12'd2684: out <= 24'hac82d4;
        12'd2685: out <= 24'hae85e6;
        12'd2686: out <= 24'hb088f7;
        12'd2687: out <= 24'hb088f7;
        12'd2688: out <= 24'haf8f1d;
        12'd2689: out <= 24'hb1922e;
        12'd2690: out <= 24'hb39440;
        12'd2691: out <= 24'hb1924e;
        12'd2692: out <= 24'haf915b;
        12'd2693: out <= 24'hb2946c;
        12'd2694: out <= 24'hb4967e;
        12'd2695: out <= 24'hb2948b;
        12'd2696: out <= 24'hb09398;
        12'd2697: out <= 24'hb296aa;
        12'd2698: out <= 24'hb598bb;
        12'd2699: out <= 24'hb396c8;
        12'd2700: out <= 24'hb195d5;
        12'd2701: out <= 24'hb398e6;
        12'd2702: out <= 24'hb59af8;
        12'd2703: out <= 24'hb59af8;
        12'd2704: out <= 24'hb3a21e;
        12'd2705: out <= 24'hb2a02c;
        12'd2706: out <= 24'hb4a23d;
        12'd2707: out <= 24'hb6a54e;
        12'd2708: out <= 24'hb4a45c;
        12'd2709: out <= 24'hb2a26a;
        12'd2710: out <= 24'hb4a47b;
        12'd2711: out <= 24'hb6a78c;
        12'd2712: out <= 24'hb4a699;
        12'd2713: out <= 24'hb2a4a6;
        12'd2714: out <= 24'hb5a6b8;
        12'd2715: out <= 24'hb7a9ca;
        12'd2716: out <= 24'hb5a8d6;
        12'd2717: out <= 24'hb4a6e4;
        12'd2718: out <= 24'hb6a8f5;
        12'd2719: out <= 24'hb6a8f5;
        12'd2720: out <= 24'hb7b520;
        12'd2721: out <= 24'hb6b32d;
        12'd2722: out <= 24'hb4b13a;
        12'd2723: out <= 24'hb6b44c;
        12'd2724: out <= 24'hb8b65d;
        12'd2725: out <= 24'hb6b46a;
        12'd2726: out <= 24'hb4b378;
        12'd2727: out <= 24'hb6b689;
        12'd2728: out <= 24'hb9b89a;
        12'd2729: out <= 24'hb7b6a8;
        12'd2730: out <= 24'hb5b5b5;
        12'd2731: out <= 24'hb7b8c6;
        12'd2732: out <= 24'hb9bad8;
        12'd2733: out <= 24'hb8b8e5;
        12'd2734: out <= 24'hb6b7f2;
        12'd2735: out <= 24'hb6b7f2;
        12'd2736: out <= 24'hb8c41d;
        12'd2737: out <= 24'hbac62e;
        12'd2738: out <= 24'hb8c43c;
        12'd2739: out <= 24'hb6c248;
        12'd2740: out <= 24'hb8c45a;
        12'd2741: out <= 24'hbac76c;
        12'd2742: out <= 24'hb8c679;
        12'd2743: out <= 24'hb6c486;
        12'd2744: out <= 24'hb9c697;
        12'd2745: out <= 24'hbcc9a8;
        12'd2746: out <= 24'hbac8b6;
        12'd2747: out <= 24'hb8c6c4;
        12'd2748: out <= 24'hbac8d5;
        12'd2749: out <= 24'hbccbe6;
        12'd2750: out <= 24'hbacaf4;
        12'd2751: out <= 24'hbacaf4;
        12'd2752: out <= 24'hb8d21a;
        12'd2753: out <= 24'hbad42c;
        12'd2754: out <= 24'hbcd73d;
        12'd2755: out <= 24'hbad54a;
        12'd2756: out <= 24'hb9d357;
        12'd2757: out <= 24'hbbd668;
        12'd2758: out <= 24'hbdd87a;
        12'd2759: out <= 24'hbbd687;
        12'd2760: out <= 24'hb9d594;
        12'd2761: out <= 24'hbcd8a6;
        12'd2762: out <= 24'hbedab7;
        12'd2763: out <= 24'hbcd8c4;
        12'd2764: out <= 24'hbad7d2;
        12'd2765: out <= 24'hbcdae4;
        12'd2766: out <= 24'hbedcf5;
        12'd2767: out <= 24'hbedcf5;
        12'd2768: out <= 24'hbce41b;
        12'd2769: out <= 24'hbae328;
        12'd2770: out <= 24'hbce63a;
        12'd2771: out <= 24'hbee84b;
        12'd2772: out <= 24'hbde658;
        12'd2773: out <= 24'hbbe466;
        12'd2774: out <= 24'hbde677;
        12'd2775: out <= 24'hc0e988;
        12'd2776: out <= 24'hbee896;
        12'd2777: out <= 24'hbce6a2;
        12'd2778: out <= 24'hbee8b4;
        12'd2779: out <= 24'hc0ebc6;
        12'd2780: out <= 24'hbeead3;
        12'd2781: out <= 24'hbce8e0;
        12'd2782: out <= 24'hbeeaf2;
        12'd2783: out <= 24'hbeeaf2;
        12'd2784: out <= 24'hc1f71c;
        12'd2785: out <= 24'hbff62a;
        12'd2786: out <= 24'hbdf437;
        12'd2787: out <= 24'hbff648;
        12'd2788: out <= 24'hc1f959;
        12'd2789: out <= 24'hbff766;
        12'd2790: out <= 24'hbdf574;
        12'd2791: out <= 24'hc0f886;
        12'd2792: out <= 24'hc2fa97;
        12'd2793: out <= 24'hc0f8a4;
        12'd2794: out <= 24'hbef7b1;
        12'd2795: out <= 24'hc0fac2;
        12'd2796: out <= 24'hc3fcd4;
        12'd2797: out <= 24'hc1fae2;
        12'd2798: out <= 24'hbff9ef;
        12'd2799: out <= 24'hbff9ef;
        12'd2800: out <= 24'hc1f71c;
        12'd2801: out <= 24'hbff62a;
        12'd2802: out <= 24'hbdf437;
        12'd2803: out <= 24'hbff648;
        12'd2804: out <= 24'hc1f959;
        12'd2805: out <= 24'hbff766;
        12'd2806: out <= 24'hbdf574;
        12'd2807: out <= 24'hc0f886;
        12'd2808: out <= 24'hc2fa97;
        12'd2809: out <= 24'hc0f8a4;
        12'd2810: out <= 24'hbef7b1;
        12'd2811: out <= 24'hc0fac2;
        12'd2812: out <= 24'hc3fcd4;
        12'd2813: out <= 24'hc1fae2;
        12'd2814: out <= 24'hbff9ef;
        12'd2815: out <= 24'hbff9ef;
        12'd2816: out <= 24'haa0a27;
        12'd2817: out <= 24'ha80934;
        12'd2818: out <= 24'ha70842;
        12'd2819: out <= 24'ha90a52;
        12'd2820: out <= 24'hab0c64;
        12'd2821: out <= 24'ha90b72;
        12'd2822: out <= 24'ha70a7f;
        12'd2823: out <= 24'haa0c90;
        12'd2824: out <= 24'hac0ea2;
        12'd2825: out <= 24'haa0caf;
        12'd2826: out <= 24'ha80bbc;
        12'd2827: out <= 24'haa0ece;
        12'd2828: out <= 24'hac10df;
        12'd2829: out <= 24'haa0eec;
        12'd2830: out <= 24'ha90cfa;
        12'd2831: out <= 24'ha90cfa;
        12'd2832: out <= 24'hae1d28;
        12'd2833: out <= 24'hac1c36;
        12'd2834: out <= 24'hab1a42;
        12'd2835: out <= 24'hae1c54;
        12'd2836: out <= 24'hb01f66;
        12'd2837: out <= 24'hae1e72;
        12'd2838: out <= 24'hac1c80;
        12'd2839: out <= 24'hae1e92;
        12'd2840: out <= 24'hb021a3;
        12'd2841: out <= 24'hae20b0;
        12'd2842: out <= 24'hac1ebd;
        12'd2843: out <= 24'hae20ce;
        12'd2844: out <= 24'hb023e0;
        12'd2845: out <= 24'hae21ee;
        12'd2846: out <= 24'had1ffa;
        12'd2847: out <= 24'had1ffa;
        12'd2848: out <= 24'haf2c25;
        12'd2849: out <= 24'had2a32;
        12'd2850: out <= 24'haf2c44;
        12'd2851: out <= 24'hb22f56;
        12'd2852: out <= 24'hb02e62;
        12'd2853: out <= 24'hae2c70;
        12'd2854: out <= 24'hb02e81;
        12'd2855: out <= 24'hb23192;
        12'd2856: out <= 24'hb030a0;
        12'd2857: out <= 24'hae2ead;
        12'd2858: out <= 24'hb130be;
        12'd2859: out <= 24'hb333d0;
        12'd2860: out <= 24'hb131dd;
        12'd2861: out <= 24'haf2fea;
        12'd2862: out <= 24'hb132fc;
        12'd2863: out <= 24'hb132fc;
        12'd2864: out <= 24'hb03a22;
        12'd2865: out <= 24'hb23c34;
        12'd2866: out <= 24'hb43f45;
        12'd2867: out <= 24'hb23e52;
        12'd2868: out <= 24'hb03c60;
        12'd2869: out <= 24'hb23e70;
        12'd2870: out <= 24'hb44182;
        12'd2871: out <= 24'hb24090;
        12'd2872: out <= 24'hb03e9d;
        12'd2873: out <= 24'hb240ae;
        12'd2874: out <= 24'hb543c0;
        12'd2875: out <= 24'hb442cc;
        12'd2876: out <= 24'hb240da;
        12'd2877: out <= 24'hb442eb;
        12'd2878: out <= 24'hb644fc;
        12'd2879: out <= 24'hb644fc;
        12'd2880: out <= 24'hb44c23;
        12'd2881: out <= 24'hb64f34;
        12'd2882: out <= 24'hb44e42;
        12'd2883: out <= 24'hb24c50;
        12'd2884: out <= 24'hb44e61;
        12'd2885: out <= 24'hb65172;
        12'd2886: out <= 24'hb4507f;
        12'd2887: out <= 24'hb24e8c;
        12'd2888: out <= 24'hb5509e;
        12'd2889: out <= 24'hb753b0;
        12'd2890: out <= 24'hb552bc;
        12'd2891: out <= 24'hb450ca;
        12'd2892: out <= 24'hb652db;
        12'd2893: out <= 24'hb855ec;
        12'd2894: out <= 24'hb653fa;
        12'd2895: out <= 24'hb653fa;
        12'd2896: out <= 24'hb86024;
        12'd2897: out <= 24'hb65e32;
        12'd2898: out <= 24'hb45c3f;
        12'd2899: out <= 24'hb65e50;
        12'd2900: out <= 24'hb86162;
        12'd2901: out <= 24'hb6606f;
        12'd2902: out <= 24'hb45e7c;
        12'd2903: out <= 24'hb7608e;
        12'd2904: out <= 24'hba639f;
        12'd2905: out <= 24'hb862ac;
        12'd2906: out <= 24'hb660ba;
        12'd2907: out <= 24'hb862cb;
        12'd2908: out <= 24'hba65dc;
        12'd2909: out <= 24'hb864ea;
        12'd2910: out <= 24'hb662f7;
        12'd2911: out <= 24'hb662f7;
        12'd2912: out <= 24'hb86e22;
        12'd2913: out <= 24'hb66c2e;
        12'd2914: out <= 24'hb86e40;
        12'd2915: out <= 24'hba7152;
        12'd2916: out <= 24'hb9705f;
        12'd2917: out <= 24'hb76e6c;
        12'd2918: out <= 24'hb9707d;
        12'd2919: out <= 24'hbc738e;
        12'd2920: out <= 24'hba729c;
        12'd2921: out <= 24'hb870aa;
        12'd2922: out <= 24'hba72bb;
        12'd2923: out <= 24'hbc75cc;
        12'd2924: out <= 24'hba74da;
        12'd2925: out <= 24'hb872e6;
        12'd2926: out <= 24'hba74f8;
        12'd2927: out <= 24'hba74f8;
        12'd2928: out <= 24'hb87c1e;
        12'd2929: out <= 24'hba7e30;
        12'd2930: out <= 24'hbc8141;
        12'd2931: out <= 24'hba804e;
        12'd2932: out <= 24'hb97e5c;
        12'd2933: out <= 24'hbc806e;
        12'd2934: out <= 24'hbe837e;
        12'd2935: out <= 24'hbc828c;
        12'd2936: out <= 24'hba8099;
        12'd2937: out <= 24'hbc82aa;
        12'd2938: out <= 24'hbe85bc;
        12'd2939: out <= 24'hbc84ca;
        12'd2940: out <= 24'hba82d6;
        12'd2941: out <= 24'hbc84e8;
        12'd2942: out <= 24'hbe87f9;
        12'd2943: out <= 24'hbe87f9;
        12'd2944: out <= 24'hbd8e20;
        12'd2945: out <= 24'hbf9130;
        12'd2946: out <= 24'hc19442;
        12'd2947: out <= 24'hbf9250;
        12'd2948: out <= 24'hbd905d;
        12'd2949: out <= 24'hc0936e;
        12'd2950: out <= 24'hc29680;
        12'd2951: out <= 24'hc0948d;
        12'd2952: out <= 24'hbe929a;
        12'd2953: out <= 24'hc095ac;
        12'd2954: out <= 24'hc398bd;
        12'd2955: out <= 24'hc196ca;
        12'd2956: out <= 24'hbf94d8;
        12'd2957: out <= 24'hc197e8;
        12'd2958: out <= 24'hc39afa;
        12'd2959: out <= 24'hc39afa;
        12'd2960: out <= 24'hc1a220;
        12'd2961: out <= 24'hc4a432;
        12'd2962: out <= 24'hc6a644;
        12'd2963: out <= 24'hc4a450;
        12'd2964: out <= 24'hc2a35e;
        12'd2965: out <= 24'hc4a670;
        12'd2966: out <= 24'hc6a881;
        12'd2967: out <= 24'hc4a68e;
        12'd2968: out <= 24'hc2a59b;
        12'd2969: out <= 24'hc0a4a8;
        12'd2970: out <= 24'hc3a6ba;
        12'd2971: out <= 24'hc5a8cc;
        12'd2972: out <= 24'hc3a7d8;
        12'd2973: out <= 24'hc2a6e6;
        12'd2974: out <= 24'hc4a8f7;
        12'd2975: out <= 24'hc4a8f7;
        12'd2976: out <= 24'hc5b422;
        12'd2977: out <= 24'hc8b734;
        12'd2978: out <= 24'hc6b540;
        12'd2979: out <= 24'hc4b34e;
        12'd2980: out <= 24'hc6b65f;
        12'd2981: out <= 24'hc8b870;
        12'd2982: out <= 24'hc6b67e;
        12'd2983: out <= 24'hc4b58b;
        12'd2984: out <= 24'hc7b89c;
        12'd2985: out <= 24'hc5b6aa;
        12'd2986: out <= 24'hc3b4b7;
        12'd2987: out <= 24'hc5b7c8;
        12'd2988: out <= 24'hc7bada;
        12'd2989: out <= 24'hc6b8e7;
        12'd2990: out <= 24'hc4b6f4;
        12'd2991: out <= 24'hc4b6f4;
        12'd2992: out <= 24'hcac723;
        12'd2993: out <= 24'hc8c630;
        12'd2994: out <= 24'hc6c43e;
        12'd2995: out <= 24'hc8c64e;
        12'd2996: out <= 24'hcac860;
        12'd2997: out <= 24'hc8c66e;
        12'd2998: out <= 24'hc6c57b;
        12'd2999: out <= 24'hc8c88c;
        12'd3000: out <= 24'hcbca9e;
        12'd3001: out <= 24'hcac8aa;
        12'd3002: out <= 24'hc8c7b8;
        12'd3003: out <= 24'hcacaca;
        12'd3004: out <= 24'hccccdb;
        12'd3005: out <= 24'hcacae8;
        12'd3006: out <= 24'hc8c9f6;
        12'd3007: out <= 24'hc8c9f6;
        12'd3008: out <= 24'hcad620;
        12'd3009: out <= 24'hc8d42e;
        12'd3010: out <= 24'hcad63f;
        12'd3011: out <= 24'hccd950;
        12'd3012: out <= 24'hcbd75d;
        12'd3013: out <= 24'hc9d56a;
        12'd3014: out <= 24'hcbd87c;
        12'd3015: out <= 24'hcdda8e;
        12'd3016: out <= 24'hcbd89a;
        12'd3017: out <= 24'hcad7a8;
        12'd3018: out <= 24'hccdab9;
        12'd3019: out <= 24'hcedcca;
        12'd3020: out <= 24'hccdad8;
        12'd3021: out <= 24'hcad9e6;
        12'd3022: out <= 24'hccdcf7;
        12'd3023: out <= 24'hccdcf7;
        12'd3024: out <= 24'hcae41d;
        12'd3025: out <= 24'hcce62e;
        12'd3026: out <= 24'hcee940;
        12'd3027: out <= 24'hcce84d;
        12'd3028: out <= 24'hcbe65a;
        12'd3029: out <= 24'hcee86c;
        12'd3030: out <= 24'hd0ea7d;
        12'd3031: out <= 24'hcee88a;
        12'd3032: out <= 24'hcce798;
        12'd3033: out <= 24'hceeaa9;
        12'd3034: out <= 24'hd0ecba;
        12'd3035: out <= 24'hceeac8;
        12'd3036: out <= 24'hcce9d5;
        12'd3037: out <= 24'hceebe6;
        12'd3038: out <= 24'hd0eef8;
        12'd3039: out <= 24'hd0eef8;
        12'd3040: out <= 24'hcff61e;
        12'd3041: out <= 24'hd1f930;
        12'd3042: out <= 24'hcff83d;
        12'd3043: out <= 24'hcdf64a;
        12'd3044: out <= 24'hcff85b;
        12'd3045: out <= 24'hd2fb6c;
        12'd3046: out <= 24'hd0f97a;
        12'd3047: out <= 24'hcef788;
        12'd3048: out <= 24'hd0fa99;
        12'd3049: out <= 24'hd2fcaa;
        12'd3050: out <= 24'hd0fab8;
        12'd3051: out <= 24'hcef9c4;
        12'd3052: out <= 24'hd1fcd6;
        12'd3053: out <= 24'hd3fee8;
        12'd3054: out <= 24'hd1fcf5;
        12'd3055: out <= 24'hd1fcf5;
        12'd3056: out <= 24'hcff61e;
        12'd3057: out <= 24'hd1f930;
        12'd3058: out <= 24'hcff83d;
        12'd3059: out <= 24'hcdf64a;
        12'd3060: out <= 24'hcff85b;
        12'd3061: out <= 24'hd2fb6c;
        12'd3062: out <= 24'hd0f97a;
        12'd3063: out <= 24'hcef788;
        12'd3064: out <= 24'hd0fa99;
        12'd3065: out <= 24'hd2fcaa;
        12'd3066: out <= 24'hd0fab8;
        12'd3067: out <= 24'hcef9c4;
        12'd3068: out <= 24'hd1fcd6;
        12'd3069: out <= 24'hd3fee8;
        12'd3070: out <= 24'hd1fcf5;
        12'd3071: out <= 24'hd1fcf5;
        12'd3072: out <= 24'hb80a29;
        12'd3073: out <= 24'hb60836;
        12'd3074: out <= 24'hb50744;
        12'd3075: out <= 24'hb70a55;
        12'd3076: out <= 24'hb90c66;
        12'd3077: out <= 24'hb70a74;
        12'd3078: out <= 24'hb50981;
        12'd3079: out <= 24'hb80c92;
        12'd3080: out <= 24'hba0ea4;
        12'd3081: out <= 24'hb80cb1;
        12'd3082: out <= 24'hb60abe;
        12'd3083: out <= 24'hb80cd0;
        12'd3084: out <= 24'hba0fe1;
        12'd3085: out <= 24'hb80eee;
        12'd3086: out <= 24'hb70cfc;
        12'd3087: out <= 24'hb70cfc;
        12'd3088: out <= 24'hbc1c2a;
        12'd3089: out <= 24'hba1b38;
        12'd3090: out <= 24'hb91a45;
        12'd3091: out <= 24'hbc1c56;
        12'd3092: out <= 24'hbe1e68;
        12'd3093: out <= 24'hbc1d74;
        12'd3094: out <= 24'hba1c82;
        12'd3095: out <= 24'hbc1e94;
        12'd3096: out <= 24'hbe20a5;
        12'd3097: out <= 24'hbc1fb2;
        12'd3098: out <= 24'hba1dbf;
        12'd3099: out <= 24'hbc20d0;
        12'd3100: out <= 24'hbe22e2;
        12'd3101: out <= 24'hbc20f0;
        12'd3102: out <= 24'hbb1efd;
        12'd3103: out <= 24'hbb1efd;
        12'd3104: out <= 24'hc12f2b;
        12'd3105: out <= 24'hbf2e38;
        12'd3106: out <= 24'hbd2c46;
        12'd3107: out <= 24'hc02e58;
        12'd3108: out <= 24'hc23169;
        12'd3109: out <= 24'hc03076;
        12'd3110: out <= 24'hbe2e83;
        12'd3111: out <= 24'hc03094;
        12'd3112: out <= 24'hc233a6;
        12'd3113: out <= 24'hc032b3;
        12'd3114: out <= 24'hbf30c0;
        12'd3115: out <= 24'hc132d2;
        12'd3116: out <= 24'hc335e3;
        12'd3117: out <= 24'hc133f0;
        12'd3118: out <= 24'hbf31fe;
        12'd3119: out <= 24'hbf31fe;
        12'd3120: out <= 24'hc23e28;
        12'd3121: out <= 24'hc4403a;
        12'd3122: out <= 24'hc23e47;
        12'd3123: out <= 24'hc03d54;
        12'd3124: out <= 24'hc24066;
        12'd3125: out <= 24'hc44277;
        12'd3126: out <= 24'hc24084;
        12'd3127: out <= 24'hc03f92;
        12'd3128: out <= 24'hc242a3;
        12'd3129: out <= 24'hc444b4;
        12'd3130: out <= 24'hc342c2;
        12'd3131: out <= 24'hc241ce;
        12'd3132: out <= 24'hc444e0;
        12'd3133: out <= 24'hc646f1;
        12'd3134: out <= 24'hc444fe;
        12'd3135: out <= 24'hc444fe;
        12'd3136: out <= 24'hc24c25;
        12'd3137: out <= 24'hc44e36;
        12'd3138: out <= 24'hc65148;
        12'd3139: out <= 24'hc45056;
        12'd3140: out <= 24'hc24e63;
        12'd3141: out <= 24'hc45074;
        12'd3142: out <= 24'hc75385;
        12'd3143: out <= 24'hc55292;
        12'd3144: out <= 24'hc350a0;
        12'd3145: out <= 24'hc552b2;
        12'd3146: out <= 24'hc755c3;
        12'd3147: out <= 24'hc654d0;
        12'd3148: out <= 24'hc452dd;
        12'd3149: out <= 24'hc654ee;
        12'd3150: out <= 24'hc857ff;
        12'd3151: out <= 24'hc857ff;
        12'd3152: out <= 24'hc65f26;
        12'd3153: out <= 24'hc45d34;
        12'd3154: out <= 24'hc66045;
        12'd3155: out <= 24'hc86256;
        12'd3156: out <= 24'hc66064;
        12'd3157: out <= 24'hc45f71;
        12'd3158: out <= 24'hc76282;
        12'd3159: out <= 24'hca6494;
        12'd3160: out <= 24'hc862a1;
        12'd3161: out <= 24'hc661ae;
        12'd3162: out <= 24'hc864c0;
        12'd3163: out <= 24'hca66d2;
        12'd3164: out <= 24'hc864de;
        12'd3165: out <= 24'hc663ec;
        12'd3166: out <= 24'hc866fc;
        12'd3167: out <= 24'hc866fc;
        12'd3168: out <= 24'hca7228;
        12'd3169: out <= 24'hc87035;
        12'd3170: out <= 24'hc66e42;
        12'd3171: out <= 24'hc87054;
        12'd3172: out <= 24'hcb7365;
        12'd3173: out <= 24'hc97272;
        12'd3174: out <= 24'hc7707f;
        12'd3175: out <= 24'hca7290;
        12'd3176: out <= 24'hcc75a2;
        12'd3177: out <= 24'hca74b0;
        12'd3178: out <= 24'hc872bd;
        12'd3179: out <= 24'hca74ce;
        12'd3180: out <= 24'hcc77e0;
        12'd3181: out <= 24'hca76ed;
        12'd3182: out <= 24'hc874fa;
        12'd3183: out <= 24'hc874fa;
        12'd3184: out <= 24'hca8025;
        12'd3185: out <= 24'hcc8236;
        12'd3186: out <= 24'hca8043;
        12'd3187: out <= 24'hc87f50;
        12'd3188: out <= 24'hcb8262;
        12'd3189: out <= 24'hce8474;
        12'd3190: out <= 24'hcc8280;
        12'd3191: out <= 24'hca818e;
        12'd3192: out <= 24'hcc849f;
        12'd3193: out <= 24'hce86b0;
        12'd3194: out <= 24'hcc84be;
        12'd3195: out <= 24'hca83cc;
        12'd3196: out <= 24'hcc86dd;
        12'd3197: out <= 24'hce88ee;
        12'd3198: out <= 24'hcc86fb;
        12'd3199: out <= 24'hcc86fb;
        12'd3200: out <= 24'hcb8e22;
        12'd3201: out <= 24'hcd9033;
        12'd3202: out <= 24'hcf9344;
        12'd3203: out <= 24'hcd9252;
        12'd3204: out <= 24'hcb905f;
        12'd3205: out <= 24'hce9270;
        12'd3206: out <= 24'hd09582;
        12'd3207: out <= 24'hce948f;
        12'd3208: out <= 24'hcc929c;
        12'd3209: out <= 24'hce94ae;
        12'd3210: out <= 24'hd197bf;
        12'd3211: out <= 24'hcf96cc;
        12'd3212: out <= 24'hcd94da;
        12'd3213: out <= 24'hcf96eb;
        12'd3214: out <= 24'hd199fc;
        12'd3215: out <= 24'hd199fc;
        12'd3216: out <= 24'hcfa123;
        12'd3217: out <= 24'hd2a434;
        12'd3218: out <= 24'hd4a646;
        12'd3219: out <= 24'hd2a452;
        12'd3220: out <= 24'hd0a260;
        12'd3221: out <= 24'hd2a572;
        12'd3222: out <= 24'hd4a883;
        12'd3223: out <= 24'hd2a690;
        12'd3224: out <= 24'hd0a49d;
        12'd3225: out <= 24'hcea3aa;
        12'd3226: out <= 24'hd1a6bc;
        12'd3227: out <= 24'hd3a8ce;
        12'd3228: out <= 24'hd1a6db;
        12'd3229: out <= 24'hd0a5e8;
        12'd3230: out <= 24'hd2a8f9;
        12'd3231: out <= 24'hd2a8f9;
        12'd3232: out <= 24'hd3b424;
        12'd3233: out <= 24'hd6b636;
        12'd3234: out <= 24'hd8b947;
        12'd3235: out <= 24'hd6b754;
        12'd3236: out <= 24'hd4b561;
        12'd3237: out <= 24'hd6b872;
        12'd3238: out <= 24'hd9ba84;
        12'd3239: out <= 24'hd7b891;
        12'd3240: out <= 24'hd5b79e;
        12'd3241: out <= 24'hd3b6ac;
        12'd3242: out <= 24'hd1b4b9;
        12'd3243: out <= 24'hd3b6ca;
        12'd3244: out <= 24'hd5b9dc;
        12'd3245: out <= 24'hd4b8e9;
        12'd3246: out <= 24'hd2b6f6;
        12'd3247: out <= 24'hd2b6f6;
        12'd3248: out <= 24'hd8c625;
        12'd3249: out <= 24'hd6c532;
        12'd3250: out <= 24'hd8c844;
        12'd3251: out <= 24'hdaca55;
        12'd3252: out <= 24'hd8c862;
        12'd3253: out <= 24'hd6c670;
        12'd3254: out <= 24'hd9c881;
        12'd3255: out <= 24'hdbcb92;
        12'd3256: out <= 24'hd9caa0;
        12'd3257: out <= 24'hd8c8ac;
        12'd3258: out <= 24'hd6c6ba;
        12'd3259: out <= 24'hd8c9cc;
        12'd3260: out <= 24'hdaccdd;
        12'd3261: out <= 24'hd8caea;
        12'd3262: out <= 24'hd6c8f8;
        12'd3263: out <= 24'hd6c8f8;
        12'd3264: out <= 24'hdcd926;
        12'd3265: out <= 24'hdad834;
        12'd3266: out <= 24'hd8d641;
        12'd3267: out <= 24'hdad852;
        12'd3268: out <= 24'hdddb63;
        12'd3269: out <= 24'hdbd970;
        12'd3270: out <= 24'hd9d77e;
        12'd3271: out <= 24'hdbda90;
        12'd3272: out <= 24'hdddca1;
        12'd3273: out <= 24'hdcdaae;
        12'd3274: out <= 24'hdad9bb;
        12'd3275: out <= 24'hdcdccc;
        12'd3276: out <= 24'hdedede;
        12'd3277: out <= 24'hdcdcec;
        12'd3278: out <= 24'hdadbf9;
        12'd3279: out <= 24'hdadbf9;
        12'd3280: out <= 24'hdce823;
        12'd3281: out <= 24'hdeea34;
        12'd3282: out <= 24'hdce842;
        12'd3283: out <= 24'hdae74f;
        12'd3284: out <= 24'hddea60;
        12'd3285: out <= 24'he0ec72;
        12'd3286: out <= 24'hdeea7f;
        12'd3287: out <= 24'hdce88c;
        12'd3288: out <= 24'hdeea9e;
        12'd3289: out <= 24'he0edb0;
        12'd3290: out <= 24'hdeecbc;
        12'd3291: out <= 24'hdceaca;
        12'd3292: out <= 24'hdeecdb;
        12'd3293: out <= 24'he0eeec;
        12'd3294: out <= 24'hdeedfa;
        12'd3295: out <= 24'hdeedfa;
        12'd3296: out <= 24'hddf620;
        12'd3297: out <= 24'hdff832;
        12'd3298: out <= 24'he1fb43;
        12'd3299: out <= 24'hdffa50;
        12'd3300: out <= 24'hddf85d;
        12'd3301: out <= 24'he0fa6e;
        12'd3302: out <= 24'he2fd80;
        12'd3303: out <= 24'he0fb8e;
        12'd3304: out <= 24'hdef99b;
        12'd3305: out <= 24'he0fcac;
        12'd3306: out <= 24'he2febe;
        12'd3307: out <= 24'he0fccb;
        12'd3308: out <= 24'hdffbd8;
        12'd3309: out <= 24'he1fdea;
        12'd3310: out <= 24'he3fffb;
        12'd3311: out <= 24'he3fffb;
        12'd3312: out <= 24'hddf620;
        12'd3313: out <= 24'hdff832;
        12'd3314: out <= 24'he1fb43;
        12'd3315: out <= 24'hdffa50;
        12'd3316: out <= 24'hddf85d;
        12'd3317: out <= 24'he0fa6e;
        12'd3318: out <= 24'he2fd80;
        12'd3319: out <= 24'he0fb8e;
        12'd3320: out <= 24'hdef99b;
        12'd3321: out <= 24'he0fcac;
        12'd3322: out <= 24'he2febe;
        12'd3323: out <= 24'he0fccb;
        12'd3324: out <= 24'hdffbd8;
        12'd3325: out <= 24'he1fdea;
        12'd3326: out <= 24'he3fffb;
        12'd3327: out <= 24'he3fffb;
        12'd3328: out <= 24'hc60a2b;
        12'd3329: out <= 24'hc80c3c;
        12'd3330: out <= 24'hc70a4a;
        12'd3331: out <= 24'hc50957;
        12'd3332: out <= 24'hc70c68;
        12'd3333: out <= 24'hca0e7a;
        12'd3334: out <= 24'hc80c87;
        12'd3335: out <= 24'hc60b94;
        12'd3336: out <= 24'hc80ea6;
        12'd3337: out <= 24'hca10b8;
        12'd3338: out <= 24'hc80ec4;
        12'd3339: out <= 24'hc60cd2;
        12'd3340: out <= 24'hc80ee3;
        12'd3341: out <= 24'hca11f0;
        12'd3342: out <= 24'hc910fe;
        12'd3343: out <= 24'hc910fe;
        12'd3344: out <= 24'hca1c2c;
        12'd3345: out <= 24'hc81a3a;
        12'd3346: out <= 24'hc71947;
        12'd3347: out <= 24'hca1c58;
        12'd3348: out <= 24'hcc1e6a;
        12'd3349: out <= 24'hca1c76;
        12'd3350: out <= 24'hc81b84;
        12'd3351: out <= 24'hca1e96;
        12'd3352: out <= 24'hcc20a7;
        12'd3353: out <= 24'hca1eb4;
        12'd3354: out <= 24'hc81cc2;
        12'd3355: out <= 24'hca1fd2;
        12'd3356: out <= 24'hcc22e4;
        12'd3357: out <= 24'hca20f0;
        12'd3358: out <= 24'hc91efe;
        12'd3359: out <= 24'hc91efe;
        12'd3360: out <= 24'hcf2e2d;
        12'd3361: out <= 24'hcd2d3a;
        12'd3362: out <= 24'hcb2c48;
        12'd3363: out <= 24'hce2e5a;
        12'd3364: out <= 24'hd0306b;
        12'd3365: out <= 24'hce2f78;
        12'd3366: out <= 24'hcc2e85;
        12'd3367: out <= 24'hce3096;
        12'd3368: out <= 24'hd032a8;
        12'd3369: out <= 24'hce31b6;
        12'd3370: out <= 24'hcd30c2;
        12'd3371: out <= 24'hcf32d4;
        12'd3372: out <= 24'hd134e5;
        12'd3373: out <= 24'hcf32f1;
        12'd3374: out <= 24'hcd30fe;
        12'd3375: out <= 24'hcd30fe;
        12'd3376: out <= 24'hd4422e;
        12'd3377: out <= 24'hd2403c;
        12'd3378: out <= 24'hd03e49;
        12'd3379: out <= 24'hd2405a;
        12'd3380: out <= 24'hd4436c;
        12'd3381: out <= 24'hd24279;
        12'd3382: out <= 24'hd04086;
        12'd3383: out <= 24'hce3e94;
        12'd3384: out <= 24'hd041a5;
        12'd3385: out <= 24'hd244b6;
        12'd3386: out <= 24'hd142c4;
        12'd3387: out <= 24'hd040d0;
        12'd3388: out <= 24'hd243e2;
        12'd3389: out <= 24'hd446f1;
        12'd3390: out <= 24'hd244fe;
        12'd3391: out <= 24'hd244fe;
        12'd3392: out <= 24'hd4502c;
        12'd3393: out <= 24'hd24e38;
        12'd3394: out <= 24'hd4504a;
        12'd3395: out <= 24'hd6535c;
        12'd3396: out <= 24'hd45269;
        12'd3397: out <= 24'hd25076;
        12'd3398: out <= 24'hd55287;
        12'd3399: out <= 24'hd35194;
        12'd3400: out <= 24'hd150a2;
        12'd3401: out <= 24'hd352b4;
        12'd3402: out <= 24'hd554c5;
        12'd3403: out <= 24'hd453d2;
        12'd3404: out <= 24'hd252df;
        12'd3405: out <= 24'hd454ee;
        12'd3406: out <= 24'hd656ff;
        12'd3407: out <= 24'hd656ff;
        12'd3408: out <= 24'hd45e28;
        12'd3409: out <= 24'hd6603a;
        12'd3410: out <= 24'hd8634b;
        12'd3411: out <= 24'hd66258;
        12'd3412: out <= 24'hd46066;
        12'd3413: out <= 24'hd66278;
        12'd3414: out <= 24'hd96588;
        12'd3415: out <= 24'hd86496;
        12'd3416: out <= 24'hd662a3;
        12'd3417: out <= 24'hd864b4;
        12'd3418: out <= 24'hda67c6;
        12'd3419: out <= 24'hd866d4;
        12'd3420: out <= 24'hd664e0;
        12'd3421: out <= 24'hd866ee;
        12'd3422: out <= 24'hda69ff;
        12'd3423: out <= 24'hda69ff;
        12'd3424: out <= 24'hd8712a;
        12'd3425: out <= 24'hda743b;
        12'd3426: out <= 24'hd87248;
        12'd3427: out <= 24'hd67056;
        12'd3428: out <= 24'hd97267;
        12'd3429: out <= 24'hdb7578;
        12'd3430: out <= 24'hd97486;
        12'd3431: out <= 24'hd87292;
        12'd3432: out <= 24'hda74a4;
        12'd3433: out <= 24'hdc77b6;
        12'd3434: out <= 24'hda76c3;
        12'd3435: out <= 24'hd874d0;
        12'd3436: out <= 24'hda76e2;
        12'd3437: out <= 24'hdc79f0;
        12'd3438: out <= 24'hda78fc;
        12'd3439: out <= 24'hda78fc;
        12'd3440: out <= 24'hdc842b;
        12'd3441: out <= 24'hda8238;
        12'd3442: out <= 24'hd88045;
        12'd3443: out <= 24'hdb8256;
        12'd3444: out <= 24'hde8568;
        12'd3445: out <= 24'hdc8476;
        12'd3446: out <= 24'hda8282;
        12'd3447: out <= 24'hdc8494;
        12'd3448: out <= 24'hde87a6;
        12'd3449: out <= 24'hdc86b2;
        12'd3450: out <= 24'hda84c0;
        12'd3451: out <= 24'hdc86d2;
        12'd3452: out <= 24'hde89e3;
        12'd3453: out <= 24'hdc88f0;
        12'd3454: out <= 24'hda86fc;
        12'd3455: out <= 24'hda86fc;
        12'd3456: out <= 24'hdd9228;
        12'd3457: out <= 24'hdb9035;
        12'd3458: out <= 24'hdd9246;
        12'd3459: out <= 24'he09558;
        12'd3460: out <= 24'hde9465;
        12'd3461: out <= 24'hdc9272;
        12'd3462: out <= 24'hde9484;
        12'd3463: out <= 24'he09796;
        12'd3464: out <= 24'hde96a2;
        12'd3465: out <= 24'hdc94b0;
        12'd3466: out <= 24'hdf96c1;
        12'd3467: out <= 24'he199d2;
        12'd3468: out <= 24'hdf98e0;
        12'd3469: out <= 24'hdd96ec;
        12'd3470: out <= 24'hdf98fe;
        12'd3471: out <= 24'hdf98fe;
        12'd3472: out <= 24'hdda025;
        12'd3473: out <= 24'he0a336;
        12'd3474: out <= 24'he2a648;
        12'd3475: out <= 24'he0a454;
        12'd3476: out <= 24'hdea262;
        12'd3477: out <= 24'he0a474;
        12'd3478: out <= 24'he2a785;
        12'd3479: out <= 24'he0a692;
        12'd3480: out <= 24'hdea4a0;
        12'd3481: out <= 24'he0a6b0;
        12'd3482: out <= 24'he3a9c2;
        12'd3483: out <= 24'he1a8d0;
        12'd3484: out <= 24'hdfa6dd;
        12'd3485: out <= 24'he2a8ec;
        12'd3486: out <= 24'he4abfe;
        12'd3487: out <= 24'he4abfe;
        12'd3488: out <= 24'he1b426;
        12'd3489: out <= 24'he4b638;
        12'd3490: out <= 24'he6b849;
        12'd3491: out <= 24'he4b656;
        12'd3492: out <= 24'he2b463;
        12'd3493: out <= 24'he4b774;
        12'd3494: out <= 24'he7ba86;
        12'd3495: out <= 24'he5b894;
        12'd3496: out <= 24'he3b6a0;
        12'd3497: out <= 24'he5b9b2;
        12'd3498: out <= 24'he3b8bf;
        12'd3499: out <= 24'he1b6cc;
        12'd3500: out <= 24'he3b8de;
        12'd3501: out <= 24'he6bbee;
        12'd3502: out <= 24'he4bafa;
        12'd3503: out <= 24'he4bafa;
        12'd3504: out <= 24'he6c627;
        12'd3505: out <= 24'he4c434;
        12'd3506: out <= 24'he6c746;
        12'd3507: out <= 24'he8ca57;
        12'd3508: out <= 24'he6c864;
        12'd3509: out <= 24'he4c672;
        12'd3510: out <= 24'he7c883;
        12'd3511: out <= 24'he9ca94;
        12'd3512: out <= 24'he7c9a2;
        12'd3513: out <= 24'he6c8ae;
        12'd3514: out <= 24'he4c6bc;
        12'd3515: out <= 24'he6c8ce;
        12'd3516: out <= 24'he8cbdf;
        12'd3517: out <= 24'he6caec;
        12'd3518: out <= 24'he4c8fa;
        12'd3519: out <= 24'he4c8fa;
        12'd3520: out <= 24'head828;
        12'd3521: out <= 24'he8d736;
        12'd3522: out <= 24'he6d643;
        12'd3523: out <= 24'he8d854;
        12'd3524: out <= 24'hebda65;
        12'd3525: out <= 24'he9d872;
        12'd3526: out <= 24'he7d680;
        12'd3527: out <= 24'he9d992;
        12'd3528: out <= 24'hebdca3;
        12'd3529: out <= 24'headab0;
        12'd3530: out <= 24'he8d8bd;
        12'd3531: out <= 24'headbce;
        12'd3532: out <= 24'hecdee0;
        12'd3533: out <= 24'headcee;
        12'd3534: out <= 24'he8dafb;
        12'd3535: out <= 24'he8dafb;
        12'd3536: out <= 24'heeeb29;
        12'd3537: out <= 24'hecea36;
        12'd3538: out <= 24'heae844;
        12'd3539: out <= 24'hecea56;
        12'd3540: out <= 24'heeed66;
        12'd3541: out <= 24'heeeb74;
        12'd3542: out <= 24'hece981;
        12'd3543: out <= 24'heceb92;
        12'd3544: out <= 24'heeeea4;
        12'd3545: out <= 24'heeecb2;
        12'd3546: out <= 24'hecebbe;
        12'd3547: out <= 24'hececd0;
        12'd3548: out <= 24'heeeee1;
        12'd3549: out <= 24'heeeeee;
        12'd3550: out <= 24'hecedfc;
        12'd3551: out <= 24'hecedfc;
        12'd3552: out <= 24'heefa26;
        12'd3553: out <= 24'hedf834;
        12'd3554: out <= 24'heffa45;
        12'd3555: out <= 24'hf0fd56;
        12'd3556: out <= 24'heefc64;
        12'd3557: out <= 24'heefa70;
        12'd3558: out <= 24'hf0fc82;
        12'd3559: out <= 24'hf0fe94;
        12'd3560: out <= 24'heefca1;
        12'd3561: out <= 24'heefbae;
        12'd3562: out <= 24'hf0fec0;
        12'd3563: out <= 24'hf0fed1;
        12'd3564: out <= 24'heffdde;
        12'd3565: out <= 24'heffdec;
        12'd3566: out <= 24'hf1fffd;
        12'd3567: out <= 24'hf1fffd;
        12'd3568: out <= 24'heefa26;
        12'd3569: out <= 24'hedf834;
        12'd3570: out <= 24'heffa45;
        12'd3571: out <= 24'hf0fd56;
        12'd3572: out <= 24'heefc64;
        12'd3573: out <= 24'heefa70;
        12'd3574: out <= 24'hf0fc82;
        12'd3575: out <= 24'hf0fe94;
        12'd3576: out <= 24'heefca1;
        12'd3577: out <= 24'heefbae;
        12'd3578: out <= 24'hf0fec0;
        12'd3579: out <= 24'hf0fed1;
        12'd3580: out <= 24'heffdde;
        12'd3581: out <= 24'heffdec;
        12'd3582: out <= 24'hf1fffd;
        12'd3583: out <= 24'hf1fffd;
        12'd3584: out <= 24'hd4092d;
        12'd3585: out <= 24'hd60c3e;
        12'd3586: out <= 24'hd90e50;
        12'd3587: out <= 24'hd70c5d;
        12'd3588: out <= 24'hd50b6a;
        12'd3589: out <= 24'hd80e7c;
        12'd3590: out <= 24'hda108d;
        12'd3591: out <= 24'hd80e9a;
        12'd3592: out <= 24'hd60da8;
        12'd3593: out <= 24'hd810ba;
        12'd3594: out <= 24'hda12cb;
        12'd3595: out <= 24'hd810d8;
        12'd3596: out <= 24'hd60ee5;
        12'd3597: out <= 24'hd810f2;
        12'd3598: out <= 24'hdb13ff;
        12'd3599: out <= 24'hdb13ff;
        12'd3600: out <= 24'hd81c2e;
        12'd3601: out <= 24'hd61a3c;
        12'd3602: out <= 24'hd91c4d;
        12'd3603: out <= 24'hdc1f5e;
        12'd3604: out <= 24'hda1e6c;
        12'd3605: out <= 24'hd81c78;
        12'd3606: out <= 24'hda1e8a;
        12'd3607: out <= 24'hdc219c;
        12'd3608: out <= 24'hda20a9;
        12'd3609: out <= 24'hd81eb6;
        12'd3610: out <= 24'hda20c8;
        12'd3611: out <= 24'hdc23d9;
        12'd3612: out <= 24'hda21e6;
        12'd3613: out <= 24'hd81ff2;
        12'd3614: out <= 24'hdb22ff;
        12'd3615: out <= 24'hdb22ff;
        12'd3616: out <= 24'hdd2e2f;
        12'd3617: out <= 24'hdb2c3c;
        12'd3618: out <= 24'hd92b4a;
        12'd3619: out <= 24'hdc2e5c;
        12'd3620: out <= 24'hde306d;
        12'd3621: out <= 24'hdc2e7a;
        12'd3622: out <= 24'hda2d87;
        12'd3623: out <= 24'hdc3098;
        12'd3624: out <= 24'hde32aa;
        12'd3625: out <= 24'hdc30b8;
        12'd3626: out <= 24'hdb2fc5;
        12'd3627: out <= 24'hdd32d6;
        12'd3628: out <= 24'hdf34e7;
        12'd3629: out <= 24'hdd32f3;
        12'd3630: out <= 24'hdb30ff;
        12'd3631: out <= 24'hdb30ff;
        12'd3632: out <= 24'he24130;
        12'd3633: out <= 24'he03f3e;
        12'd3634: out <= 24'hde3e4b;
        12'd3635: out <= 24'he0405c;
        12'd3636: out <= 24'he2426e;
        12'd3637: out <= 24'he0417b;
        12'd3638: out <= 24'hde4088;
        12'd3639: out <= 24'hdc3e96;
        12'd3640: out <= 24'hde40a7;
        12'd3641: out <= 24'he043b8;
        12'd3642: out <= 24'hdf42c6;
        12'd3643: out <= 24'hde40d3;
        12'd3644: out <= 24'he042e4;
        12'd3645: out <= 24'he245f3;
        12'd3646: out <= 24'he043ff;
        12'd3647: out <= 24'he043ff;
        12'd3648: out <= 24'he65432;
        12'd3649: out <= 24'he4523f;
        12'd3650: out <= 24'he2504c;
        12'd3651: out <= 24'he4525e;
        12'd3652: out <= 24'he6556f;
        12'd3653: out <= 24'he4547c;
        12'd3654: out <= 24'he35289;
        12'd3655: out <= 24'he15096;
        12'd3656: out <= 24'hdf4fa4;
        12'd3657: out <= 24'he152b6;
        12'd3658: out <= 24'he354c7;
        12'd3659: out <= 24'he252d4;
        12'd3660: out <= 24'he051e1;
        12'd3661: out <= 24'he254f0;
        12'd3662: out <= 24'he456ff;
        12'd3663: out <= 24'he456ff;
        12'd3664: out <= 24'he6622f;
        12'd3665: out <= 24'he86440;
        12'd3666: out <= 24'he6624d;
        12'd3667: out <= 24'he4615a;
        12'd3668: out <= 24'he6646c;
        12'd3669: out <= 24'he8667e;
        12'd3670: out <= 24'he7648a;
        12'd3671: out <= 24'he66398;
        12'd3672: out <= 24'he462a5;
        12'd3673: out <= 24'he664b6;
        12'd3674: out <= 24'he866c8;
        12'd3675: out <= 24'he665d6;
        12'd3676: out <= 24'he464e2;
        12'd3677: out <= 24'he666f0;
        12'd3678: out <= 24'he868ff;
        12'd3679: out <= 24'he868ff;
        12'd3680: out <= 24'he6702c;
        12'd3681: out <= 24'he8723d;
        12'd3682: out <= 24'heb754e;
        12'd3683: out <= 24'he9745c;
        12'd3684: out <= 24'he77269;
        12'd3685: out <= 24'he9747a;
        12'd3686: out <= 24'heb778c;
        12'd3687: out <= 24'hea7699;
        12'd3688: out <= 24'he874a6;
        12'd3689: out <= 24'hea76b8;
        12'd3690: out <= 24'hec79c9;
        12'd3691: out <= 24'hea78d6;
        12'd3692: out <= 24'he876e4;
        12'd3693: out <= 24'hea78f2;
        12'd3694: out <= 24'hed7bff;
        12'd3695: out <= 24'hed7bff;
        12'd3696: out <= 24'hea832d;
        12'd3697: out <= 24'he8813a;
        12'd3698: out <= 24'heb844b;
        12'd3699: out <= 24'hee865c;
        12'd3700: out <= 24'hec846a;
        12'd3701: out <= 24'hea8378;
        12'd3702: out <= 24'hec8689;
        12'd3703: out <= 24'hee889a;
        12'd3704: out <= 24'hec86a8;
        12'd3705: out <= 24'hea85b4;
        12'd3706: out <= 24'hec88c6;
        12'd3707: out <= 24'hee8ad8;
        12'd3708: out <= 24'hec88e5;
        12'd3709: out <= 24'hea87f2;
        12'd3710: out <= 24'hed8aff;
        12'd3711: out <= 24'hed8aff;
        12'd3712: out <= 24'hef962e;
        12'd3713: out <= 24'hed943b;
        12'd3714: out <= 24'heb9248;
        12'd3715: out <= 24'hee945a;
        12'd3716: out <= 24'hf0976b;
        12'd3717: out <= 24'hee9678;
        12'd3718: out <= 24'hec9486;
        12'd3719: out <= 24'hee9698;
        12'd3720: out <= 24'hf099a9;
        12'd3721: out <= 24'hee98b6;
        12'd3722: out <= 24'hed96c3;
        12'd3723: out <= 24'hef98d4;
        12'd3724: out <= 24'hf19be6;
        12'd3725: out <= 24'hef9af2;
        12'd3726: out <= 24'hed98ff;
        12'd3727: out <= 24'hed98ff;
        12'd3728: out <= 24'hefa42b;
        12'd3729: out <= 24'hf2a73c;
        12'd3730: out <= 24'hf0a54a;
        12'd3731: out <= 24'heea356;
        12'd3732: out <= 24'hf0a668;
        12'd3733: out <= 24'hf2a87a;
        12'd3734: out <= 24'hf0a687;
        12'd3735: out <= 24'heea594;
        12'd3736: out <= 24'hf0a8a6;
        12'd3737: out <= 24'hf2aab7;
        12'd3738: out <= 24'hf1a8c4;
        12'd3739: out <= 24'hefa7d2;
        12'd3740: out <= 24'hf1aae3;
        12'd3741: out <= 24'hf4acf2;
        12'd3742: out <= 24'hf2aaff;
        12'd3743: out <= 24'hf2aaff;
        12'd3744: out <= 24'hefb328;
        12'd3745: out <= 24'hf2b63a;
        12'd3746: out <= 24'hf4b84b;
        12'd3747: out <= 24'hf2b658;
        12'd3748: out <= 24'hf0b465;
        12'd3749: out <= 24'hf2b676;
        12'd3750: out <= 24'hf5b988;
        12'd3751: out <= 24'hf3b896;
        12'd3752: out <= 24'hf1b6a3;
        12'd3753: out <= 24'hf3b8b4;
        12'd3754: out <= 24'hf5bbc5;
        12'd3755: out <= 24'hf3bad2;
        12'd3756: out <= 24'hf1b8e0;
        12'd3757: out <= 24'hf4baf0;
        12'd3758: out <= 24'hf6bdff;
        12'd3759: out <= 24'hf6bdff;
        12'd3760: out <= 24'hf4c629;
        12'd3761: out <= 24'hf2c436;
        12'd3762: out <= 24'hf4c648;
        12'd3763: out <= 24'hf6c959;
        12'd3764: out <= 24'hf4c766;
        12'd3765: out <= 24'hf2c574;
        12'd3766: out <= 24'hf5c885;
        12'd3767: out <= 24'hf7ca96;
        12'd3768: out <= 24'hf5c8a4;
        12'd3769: out <= 24'hf4c7b1;
        12'd3770: out <= 24'hf6cac2;
        12'd3771: out <= 24'hf8ccd4;
        12'd3772: out <= 24'hf6cae1;
        12'd3773: out <= 24'hf4c9ee;
        12'd3774: out <= 24'hf6ccfe;
        12'd3775: out <= 24'hf6ccfe;
        12'd3776: out <= 24'hf8d82a;
        12'd3777: out <= 24'hf6d638;
        12'd3778: out <= 24'hf4d545;
        12'd3779: out <= 24'hf6d856;
        12'd3780: out <= 24'hf9da67;
        12'd3781: out <= 24'hf7d874;
        12'd3782: out <= 24'hf5d682;
        12'd3783: out <= 24'hf7d894;
        12'd3784: out <= 24'hf9dba5;
        12'd3785: out <= 24'hf8dab2;
        12'd3786: out <= 24'hf6d8bf;
        12'd3787: out <= 24'hf8dad0;
        12'd3788: out <= 24'hfadde2;
        12'd3789: out <= 24'hf8dcf0;
        12'd3790: out <= 24'hf6dafd;
        12'd3791: out <= 24'hf6dafd;
        12'd3792: out <= 24'hfcea2b;
        12'd3793: out <= 24'hfae938;
        12'd3794: out <= 24'hf8e846;
        12'd3795: out <= 24'hfaea58;
        12'd3796: out <= 24'hfcec68;
        12'd3797: out <= 24'hfcea76;
        12'd3798: out <= 24'hfae883;
        12'd3799: out <= 24'hfaea94;
        12'd3800: out <= 24'hfceda6;
        12'd3801: out <= 24'hfcecb4;
        12'd3802: out <= 24'hfaeac0;
        12'd3803: out <= 24'hfaecd2;
        12'd3804: out <= 24'hfceee3;
        12'd3805: out <= 24'hfceef0;
        12'd3806: out <= 24'hfaecfe;
        12'd3807: out <= 24'hfaecfe;
        12'd3808: out <= 24'hfffd2c;
        12'd3809: out <= 24'hfefc3a;
        12'd3810: out <= 24'hfdfa47;
        12'd3811: out <= 24'hfefc58;
        12'd3812: out <= 24'hffff6a;
        12'd3813: out <= 24'hfefd77;
        12'd3814: out <= 24'hfefb84;
        12'd3815: out <= 24'hfefd96;
        12'd3816: out <= 24'hffffa7;
        12'd3817: out <= 24'hfefeb4;
        12'd3818: out <= 24'hfefdc2;
        12'd3819: out <= 24'hfefed3;
        12'd3820: out <= 24'hffffe4;
        12'd3821: out <= 24'hfffff2;
        12'd3822: out <= 24'hffffff;
        12'd3823: out <= 24'hffffff;
        12'd3824: out <= 24'hfffd2c;
        12'd3825: out <= 24'hfefc3a;
        12'd3826: out <= 24'hfdfa47;
        12'd3827: out <= 24'hfefc58;
        12'd3828: out <= 24'hffff6a;
        12'd3829: out <= 24'hfefd77;
        12'd3830: out <= 24'hfefb84;
        12'd3831: out <= 24'hfefd96;
        12'd3832: out <= 24'hffffa7;
        12'd3833: out <= 24'hfefeb4;
        12'd3834: out <= 24'hfefdc2;
        12'd3835: out <= 24'hfefed3;
        12'd3836: out <= 24'hffffe4;
        12'd3837: out <= 24'hfffff2;
        12'd3838: out <= 24'hffffff;
        12'd3839: out <= 24'hffffff;
        12'd3840: out <= 24'hd4092d;
        12'd3841: out <= 24'hd60c3e;
        12'd3842: out <= 24'hd90e50;
        12'd3843: out <= 24'hd70c5d;
        12'd3844: out <= 24'hd50b6a;
        12'd3845: out <= 24'hd80e7c;
        12'd3846: out <= 24'hda108d;
        12'd3847: out <= 24'hd80e9a;
        12'd3848: out <= 24'hd60da8;
        12'd3849: out <= 24'hd810ba;
        12'd3850: out <= 24'hda12cb;
        12'd3851: out <= 24'hd810d8;
        12'd3852: out <= 24'hd60ee5;
        12'd3853: out <= 24'hd810f2;
        12'd3854: out <= 24'hdb13ff;
        12'd3855: out <= 24'hdb13ff;
        12'd3856: out <= 24'hd81c2e;
        12'd3857: out <= 24'hd61a3c;
        12'd3858: out <= 24'hd91c4d;
        12'd3859: out <= 24'hdc1f5e;
        12'd3860: out <= 24'hda1e6c;
        12'd3861: out <= 24'hd81c78;
        12'd3862: out <= 24'hda1e8a;
        12'd3863: out <= 24'hdc219c;
        12'd3864: out <= 24'hda20a9;
        12'd3865: out <= 24'hd81eb6;
        12'd3866: out <= 24'hda20c8;
        12'd3867: out <= 24'hdc23d9;
        12'd3868: out <= 24'hda21e6;
        12'd3869: out <= 24'hd81ff2;
        12'd3870: out <= 24'hdb22ff;
        12'd3871: out <= 24'hdb22ff;
        12'd3872: out <= 24'hdd2e2f;
        12'd3873: out <= 24'hdb2c3c;
        12'd3874: out <= 24'hd92b4a;
        12'd3875: out <= 24'hdc2e5c;
        12'd3876: out <= 24'hde306d;
        12'd3877: out <= 24'hdc2e7a;
        12'd3878: out <= 24'hda2d87;
        12'd3879: out <= 24'hdc3098;
        12'd3880: out <= 24'hde32aa;
        12'd3881: out <= 24'hdc30b8;
        12'd3882: out <= 24'hdb2fc5;
        12'd3883: out <= 24'hdd32d6;
        12'd3884: out <= 24'hdf34e7;
        12'd3885: out <= 24'hdd32f3;
        12'd3886: out <= 24'hdb30ff;
        12'd3887: out <= 24'hdb30ff;
        12'd3888: out <= 24'he24130;
        12'd3889: out <= 24'he03f3e;
        12'd3890: out <= 24'hde3e4b;
        12'd3891: out <= 24'he0405c;
        12'd3892: out <= 24'he2426e;
        12'd3893: out <= 24'he0417b;
        12'd3894: out <= 24'hde4088;
        12'd3895: out <= 24'hdc3e96;
        12'd3896: out <= 24'hde40a7;
        12'd3897: out <= 24'he043b8;
        12'd3898: out <= 24'hdf42c6;
        12'd3899: out <= 24'hde40d3;
        12'd3900: out <= 24'he042e4;
        12'd3901: out <= 24'he245f3;
        12'd3902: out <= 24'he043ff;
        12'd3903: out <= 24'he043ff;
        12'd3904: out <= 24'he65432;
        12'd3905: out <= 24'he4523f;
        12'd3906: out <= 24'he2504c;
        12'd3907: out <= 24'he4525e;
        12'd3908: out <= 24'he6556f;
        12'd3909: out <= 24'he4547c;
        12'd3910: out <= 24'he35289;
        12'd3911: out <= 24'he15096;
        12'd3912: out <= 24'hdf4fa4;
        12'd3913: out <= 24'he152b6;
        12'd3914: out <= 24'he354c7;
        12'd3915: out <= 24'he252d4;
        12'd3916: out <= 24'he051e1;
        12'd3917: out <= 24'he254f0;
        12'd3918: out <= 24'he456ff;
        12'd3919: out <= 24'he456ff;
        12'd3920: out <= 24'he6622f;
        12'd3921: out <= 24'he86440;
        12'd3922: out <= 24'he6624d;
        12'd3923: out <= 24'he4615a;
        12'd3924: out <= 24'he6646c;
        12'd3925: out <= 24'he8667e;
        12'd3926: out <= 24'he7648a;
        12'd3927: out <= 24'he66398;
        12'd3928: out <= 24'he462a5;
        12'd3929: out <= 24'he664b6;
        12'd3930: out <= 24'he866c8;
        12'd3931: out <= 24'he665d6;
        12'd3932: out <= 24'he464e2;
        12'd3933: out <= 24'he666f0;
        12'd3934: out <= 24'he868ff;
        12'd3935: out <= 24'he868ff;
        12'd3936: out <= 24'he6702c;
        12'd3937: out <= 24'he8723d;
        12'd3938: out <= 24'heb754e;
        12'd3939: out <= 24'he9745c;
        12'd3940: out <= 24'he77269;
        12'd3941: out <= 24'he9747a;
        12'd3942: out <= 24'heb778c;
        12'd3943: out <= 24'hea7699;
        12'd3944: out <= 24'he874a6;
        12'd3945: out <= 24'hea76b8;
        12'd3946: out <= 24'hec79c9;
        12'd3947: out <= 24'hea78d6;
        12'd3948: out <= 24'he876e4;
        12'd3949: out <= 24'hea78f2;
        12'd3950: out <= 24'hed7bff;
        12'd3951: out <= 24'hed7bff;
        12'd3952: out <= 24'hea832d;
        12'd3953: out <= 24'he8813a;
        12'd3954: out <= 24'heb844b;
        12'd3955: out <= 24'hee865c;
        12'd3956: out <= 24'hec846a;
        12'd3957: out <= 24'hea8378;
        12'd3958: out <= 24'hec8689;
        12'd3959: out <= 24'hee889a;
        12'd3960: out <= 24'hec86a8;
        12'd3961: out <= 24'hea85b4;
        12'd3962: out <= 24'hec88c6;
        12'd3963: out <= 24'hee8ad8;
        12'd3964: out <= 24'hec88e5;
        12'd3965: out <= 24'hea87f2;
        12'd3966: out <= 24'hed8aff;
        12'd3967: out <= 24'hed8aff;
        12'd3968: out <= 24'hef962e;
        12'd3969: out <= 24'hed943b;
        12'd3970: out <= 24'heb9248;
        12'd3971: out <= 24'hee945a;
        12'd3972: out <= 24'hf0976b;
        12'd3973: out <= 24'hee9678;
        12'd3974: out <= 24'hec9486;
        12'd3975: out <= 24'hee9698;
        12'd3976: out <= 24'hf099a9;
        12'd3977: out <= 24'hee98b6;
        12'd3978: out <= 24'hed96c3;
        12'd3979: out <= 24'hef98d4;
        12'd3980: out <= 24'hf19be6;
        12'd3981: out <= 24'hef9af2;
        12'd3982: out <= 24'hed98ff;
        12'd3983: out <= 24'hed98ff;
        12'd3984: out <= 24'hefa42b;
        12'd3985: out <= 24'hf2a73c;
        12'd3986: out <= 24'hf0a54a;
        12'd3987: out <= 24'heea356;
        12'd3988: out <= 24'hf0a668;
        12'd3989: out <= 24'hf2a87a;
        12'd3990: out <= 24'hf0a687;
        12'd3991: out <= 24'heea594;
        12'd3992: out <= 24'hf0a8a6;
        12'd3993: out <= 24'hf2aab7;
        12'd3994: out <= 24'hf1a8c4;
        12'd3995: out <= 24'hefa7d2;
        12'd3996: out <= 24'hf1aae3;
        12'd3997: out <= 24'hf4acf2;
        12'd3998: out <= 24'hf2aaff;
        12'd3999: out <= 24'hf2aaff;
        12'd4000: out <= 24'hefb328;
        12'd4001: out <= 24'hf2b63a;
        12'd4002: out <= 24'hf4b84b;
        12'd4003: out <= 24'hf2b658;
        12'd4004: out <= 24'hf0b465;
        12'd4005: out <= 24'hf2b676;
        12'd4006: out <= 24'hf5b988;
        12'd4007: out <= 24'hf3b896;
        12'd4008: out <= 24'hf1b6a3;
        12'd4009: out <= 24'hf3b8b4;
        12'd4010: out <= 24'hf5bbc5;
        12'd4011: out <= 24'hf3bad2;
        12'd4012: out <= 24'hf1b8e0;
        12'd4013: out <= 24'hf4baf0;
        12'd4014: out <= 24'hf6bdff;
        12'd4015: out <= 24'hf6bdff;
        12'd4016: out <= 24'hf4c629;
        12'd4017: out <= 24'hf2c436;
        12'd4018: out <= 24'hf4c648;
        12'd4019: out <= 24'hf6c959;
        12'd4020: out <= 24'hf4c766;
        12'd4021: out <= 24'hf2c574;
        12'd4022: out <= 24'hf5c885;
        12'd4023: out <= 24'hf7ca96;
        12'd4024: out <= 24'hf5c8a4;
        12'd4025: out <= 24'hf4c7b1;
        12'd4026: out <= 24'hf6cac2;
        12'd4027: out <= 24'hf8ccd4;
        12'd4028: out <= 24'hf6cae1;
        12'd4029: out <= 24'hf4c9ee;
        12'd4030: out <= 24'hf6ccfe;
        12'd4031: out <= 24'hf6ccfe;
        12'd4032: out <= 24'hf8d82a;
        12'd4033: out <= 24'hf6d638;
        12'd4034: out <= 24'hf4d545;
        12'd4035: out <= 24'hf6d856;
        12'd4036: out <= 24'hf9da67;
        12'd4037: out <= 24'hf7d874;
        12'd4038: out <= 24'hf5d682;
        12'd4039: out <= 24'hf7d894;
        12'd4040: out <= 24'hf9dba5;
        12'd4041: out <= 24'hf8dab2;
        12'd4042: out <= 24'hf6d8bf;
        12'd4043: out <= 24'hf8dad0;
        12'd4044: out <= 24'hfadde2;
        12'd4045: out <= 24'hf8dcf0;
        12'd4046: out <= 24'hf6dafd;
        12'd4047: out <= 24'hf6dafd;
        12'd4048: out <= 24'hfcea2b;
        12'd4049: out <= 24'hfae938;
        12'd4050: out <= 24'hf8e846;
        12'd4051: out <= 24'hfaea58;
        12'd4052: out <= 24'hfcec68;
        12'd4053: out <= 24'hfcea76;
        12'd4054: out <= 24'hfae883;
        12'd4055: out <= 24'hfaea94;
        12'd4056: out <= 24'hfceda6;
        12'd4057: out <= 24'hfcecb4;
        12'd4058: out <= 24'hfaeac0;
        12'd4059: out <= 24'hfaecd2;
        12'd4060: out <= 24'hfceee3;
        12'd4061: out <= 24'hfceef0;
        12'd4062: out <= 24'hfaecfe;
        12'd4063: out <= 24'hfaecfe;
        12'd4064: out <= 24'hfffd2c;
        12'd4065: out <= 24'hfefc3a;
        12'd4066: out <= 24'hfdfa47;
        12'd4067: out <= 24'hfefc58;
        12'd4068: out <= 24'hffff6a;
        12'd4069: out <= 24'hfefd77;
        12'd4070: out <= 24'hfefb84;
        12'd4071: out <= 24'hfefd96;
        12'd4072: out <= 24'hffffa7;
        12'd4073: out <= 24'hfefeb4;
        12'd4074: out <= 24'hfefdc2;
        12'd4075: out <= 24'hfefed3;
        12'd4076: out <= 24'hffffe4;
        12'd4077: out <= 24'hfffff2;
        12'd4078: out <= 24'hffffff;
        12'd4079: out <= 24'hffffff;
        12'd4080: out <= 24'hfffd2c;
        12'd4081: out <= 24'hfefc3a;
        12'd4082: out <= 24'hfdfa47;
        12'd4083: out <= 24'hfefc58;
        12'd4084: out <= 24'hffff6a;
        12'd4085: out <= 24'hfefd77;
        12'd4086: out <= 24'hfefb84;
        12'd4087: out <= 24'hfefd96;
        12'd4088: out <= 24'hffffa7;
        12'd4089: out <= 24'hfefeb4;
        12'd4090: out <= 24'hfefdc2;
        12'd4091: out <= 24'hfefed3;
        12'd4092: out <= 24'hffffe4;
        12'd4093: out <= 24'hfffff2;
        12'd4094: out <= 24'hffffff;
        12'd4095: out <= 24'hffffff;
    endcase

endmodule
